`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/09/2022 04:08:14 AM
// Design Name: 
// Module Name: mac_array_64x64
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mac_array_64x64( clk, rst,
    ain1, ain2, ain3, ain4, ain5, ain6, ain7, ain8,
    ain9, ain10, ain11, ain12, ain13, ain14, ain15, ain16, 
    ain17, ain18, ain19, ain20, ain21, ain22, ain23, ain24, 
    ain25, ain26, ain27, ain28, ain29, ain30, ain31, ain32, 
    ain33, ain34, ain35, ain36, ain37, ain38, ain39, ain40, 
    ain41, ain42, ain43, ain44, ain45, ain46, ain47, ain48,
    ain49, ain50, ain51, ain52, ain53, ain54, ain55, ain56,
    ain57, ain58, ain59, ain60, ain61, ain62, ain63, ain64,
    
    win1, win2, win3, win4, win5, win6, win7, win8,
    win9, win10, win11, win12, win13, win14, win15, win16, 
    win17, win18, win19, win20, win21, win22, win23, win24, 
    win25, win26, win27, win28, win29, win30, win31, win32, 
    win33, win34, win35, win36, win37, win38, win39, win40, 
    win41, win42, win43, win44, win45, win46, win47, win48,
    win49, win50, win51, win52, win53, win54, win55, win56,
    win57, win58, win59, win60, win61, win62, win63, win64,
     
    sout11, sout12, sout13, sout14, sout15, sout16, sout17, sout18,
    sout19, sout1_10, sout1_11, sout1_12, sout1_13, sout1_14, sout1_15, sout1_16,
    sout1_17, sout1_18, sout1_19, sout1_20, sout1_21, sout1_22, sout1_23, sout1_24, 
    sout1_25, sout1_26, sout1_27, sout1_28, sout1_29, sout1_30, sout1_31, sout1_32,
    sout1_33, sout1_34, sout1_35, sout1_36, sout1_37, sout1_38, sout1_39, sout1_40,
    sout1_41, sout1_42, sout1_43, sout1_44, sout1_45, sout1_46, sout1_47, sout1_48,
    sout1_49, sout1_50, sout1_51, sout1_52, sout1_53, sout1_54, sout1_55, sout1_56, 
    sout1_57, sout1_58, sout1_59, sout1_60, sout1_61, sout1_62, sout1_63, sout1_64,
    
    sout21, sout22, sout23, sout24, sout25, sout26, sout27, sout28,
    sout29, sout2_10, sout2_11, sout2_12, sout2_13, sout2_14, sout2_15, sout2_16,
    sout2_17, sout2_18, sout2_19, sout2_20, sout2_21, sout2_22, sout2_23, sout2_24, 
    sout2_25, sout2_26, sout2_27, sout2_28, sout2_29, sout2_30, sout2_31, sout2_32,
    sout2_33, sout2_34, sout2_35, sout2_36, sout2_37, sout2_38, sout2_39, sout2_40,
    sout2_41, sout2_42, sout2_43, sout2_44, sout2_45, sout2_46, sout2_47, sout2_48,
    sout2_49, sout2_50, sout2_51, sout2_52, sout2_53, sout2_54, sout2_55, sout2_56, 
    sout2_57, sout2_58, sout2_59, sout2_60, sout2_61, sout2_62, sout2_63, sout2_64,
    
    sout31, sout32, sout33, sout34, sout35, sout36, sout37, sout38,
    sout39, sout3_10, sout3_11, sout3_12, sout3_13, sout3_14, sout3_15, sout3_16,
    sout3_17, sout3_18, sout3_19, sout3_20, sout3_21, sout3_22, sout3_23, sout3_24, 
    sout3_25, sout3_26, sout3_27, sout3_28, sout3_29, sout3_30, sout3_31, sout3_32,
    sout3_33, sout3_34, sout3_35, sout3_36, sout3_37, sout3_38, sout3_39, sout3_40,
    sout3_41, sout3_42, sout3_43, sout3_44, sout3_45, sout3_46, sout3_47, sout3_48,
    sout3_49, sout3_50, sout3_51, sout3_52, sout3_53, sout3_54, sout3_55, sout3_56, 
    sout3_57, sout3_58, sout3_59, sout3_60, sout3_61, sout3_62, sout3_63, sout3_64,
    
    sout41, sout42, sout43, sout44, sout45, sout46, sout47, sout48,
    sout49, sout4_10, sout4_11, sout4_12, sout4_13, sout4_14, sout4_15, sout4_16,
    sout4_17, sout4_18, sout4_19, sout4_20, sout4_21, sout4_22, sout4_23, sout4_24, 
    sout4_25, sout4_26, sout4_27, sout4_28, sout4_29, sout4_30, sout4_31, sout4_32,
    sout4_33, sout4_34, sout4_35, sout4_36, sout4_37, sout4_38, sout4_39, sout4_40,
    sout4_41, sout4_42, sout4_43, sout4_44, sout4_45, sout4_46, sout4_47, sout4_48,
    sout4_49, sout4_50, sout4_51, sout4_52, sout4_53, sout4_54, sout4_55, sout4_56, 
    sout4_57, sout4_58, sout4_59, sout4_60, sout4_61, sout4_62, sout4_63, sout4_64,
    
    sout51, sout52, sout53, sout54, sout55, sout56, sout57, sout58,
    sout59, sout5_10, sout5_11, sout5_12, sout5_13, sout5_14, sout5_15, sout5_16,
    sout5_17, sout5_18, sout5_19, sout5_20, sout5_21, sout5_22, sout5_23, sout5_24, 
    sout5_25, sout5_26, sout5_27, sout5_28, sout5_29, sout5_30, sout5_31, sout5_32,
    sout5_33, sout5_34, sout5_35, sout5_36, sout5_37, sout5_38, sout5_39, sout5_40,
    sout5_41, sout5_42, sout5_43, sout5_44, sout5_45, sout5_46, sout5_47, sout5_48,
    sout5_49, sout5_50, sout5_51, sout5_52, sout5_53, sout5_54, sout5_55, sout5_56, 
    sout5_57, sout5_58, sout5_59, sout5_60, sout5_61, sout5_62, sout5_63, sout5_64,
    
    sout61, sout62, sout63, sout64, sout65, sout66, sout67, sout68,
    sout69, sout6_10, sout6_11, sout6_12, sout6_13, sout6_14, sout6_15, sout6_16,
    sout6_17, sout6_18, sout6_19, sout6_20, sout6_21, sout6_22, sout6_23, sout6_24, 
    sout6_25, sout6_26, sout6_27, sout6_28, sout6_29, sout6_30, sout6_31, sout6_32,
    sout6_33, sout6_34, sout6_35, sout6_36, sout6_37, sout6_38, sout6_39, sout6_40,
    sout6_41, sout6_42, sout6_43, sout6_44, sout6_45, sout6_46, sout6_47, sout6_48,
    sout6_49, sout6_50, sout6_51, sout6_52, sout6_53, sout6_54, sout6_55, sout6_56, 
    sout6_57, sout6_58, sout6_59, sout6_60, sout6_61, sout6_62, sout6_63, sout6_64, 
    
    sout71, sout72, sout73, sout74, sout75, sout76, sout77, sout78,
    sout79, sout7_10, sout7_11, sout7_12, sout7_13, sout7_14, sout7_15, sout7_16,
    sout7_17, sout7_18, sout7_19, sout7_20, sout7_21, sout7_22, sout7_23, sout7_24, 
    sout7_25, sout7_26, sout7_27, sout7_28, sout7_29, sout7_30, sout7_31, sout7_32,
    sout7_33, sout7_34, sout7_35, sout7_36, sout7_37, sout7_38, sout7_39, sout7_40,
    sout7_41, sout7_42, sout7_43, sout7_44, sout7_45, sout7_46, sout7_47, sout7_48,
    sout7_49, sout7_50, sout7_51, sout7_52, sout7_53, sout7_54, sout7_55, sout7_56, 
    sout7_57, sout7_58, sout7_59, sout7_60, sout7_61, sout7_62, sout7_63, sout7_64, 
    
    sout81, sout82, sout83, sout84, sout85, sout86, sout87, sout88,
    sout89, sout8_10, sout8_11, sout8_12, sout8_13, sout8_14, sout8_15, sout8_16,
    sout8_17, sout8_18, sout8_19, sout8_20, sout8_21, sout8_22, sout8_23, sout8_24, 
    sout8_25, sout8_26, sout8_27, sout8_28, sout8_29, sout8_30, sout8_31, sout8_32,
    sout8_33, sout8_34, sout8_35, sout8_36, sout8_37, sout8_38, sout8_39, sout8_40,
    sout8_41, sout8_42, sout8_43, sout8_44, sout8_45, sout8_46, sout8_47, sout8_48,
    sout8_49, sout8_50, sout8_51, sout8_52, sout8_53, sout8_54, sout8_55, sout8_56, 
    sout8_57, sout8_58, sout8_59, sout8_60, sout8_61, sout8_62, sout8_63, sout8_64,
    
    sout91, sout92, sout93, sout94, sout95, sout96, sout97, sout98,
    sout99, sout9_10, sout9_11, sout9_12, sout9_13, sout9_14, sout9_15, sout9_16,
    sout9_17, sout9_18, sout9_19, sout9_20, sout9_21, sout9_22, sout9_23, sout9_24, 
    sout9_25, sout9_26, sout9_27, sout9_28, sout9_29, sout9_30, sout9_31, sout9_32,
    sout9_33, sout9_34, sout9_35, sout9_36, sout9_37, sout9_38, sout9_39, sout9_40,
    sout9_41, sout9_42, sout9_43, sout9_44, sout9_45, sout9_46, sout9_47, sout9_48,
    sout9_49, sout9_50, sout9_51, sout9_52, sout9_53, sout9_54, sout9_55, sout9_56, 
    sout9_57, sout9_58, sout9_59, sout9_60, sout9_61, sout9_62, sout9_63, sout9_64,
    
    sout10_1, sout10_2, sout10_3, sout10_4, sout10_5, sout10_6, sout10_7, sout10_8,
    sout10_9, sout10_10, sout10_11, sout10_12, sout10_13, sout10_14, sout10_15, sout10_16,
    sout10_17, sout10_18, sout10_19, sout10_20, sout10_21, sout10_22, sout10_23, sout10_24, 
    sout10_25, sout10_26, sout10_27, sout10_28, sout10_29, sout10_30, sout10_31, sout10_32,
    sout10_33, sout10_34, sout10_35, sout10_36, sout10_37, sout10_38, sout10_39, sout10_40,
    sout10_41, sout10_42, sout10_43, sout10_44, sout10_45, sout10_46, sout10_47, sout10_48,
    sout10_49, sout10_50, sout10_51, sout10_52, sout10_53, sout10_54, sout10_55, sout10_56, 
    sout10_57, sout10_58, sout10_59, sout10_60, sout10_61, sout10_62, sout10_63, sout10_64,
    
    sout11_1, sout11_2, sout11_3, sout11_4, sout11_5, sout11_6, sout11_7, sout11_8,
    sout11_9, sout11_10, sout11_11, sout11_12, sout11_13, sout11_14, sout11_15, sout11_16,
    sout11_17, sout11_18, sout11_19, sout11_20, sout11_21, sout11_22, sout11_23, sout11_24, 
    sout11_25, sout11_26, sout11_27, sout11_28, sout11_29, sout11_30, sout11_31, sout11_32,
    sout11_33, sout11_34, sout11_35, sout11_36, sout11_37, sout11_38, sout11_39, sout11_40,
    sout11_41, sout11_42, sout11_43, sout11_44, sout11_45, sout11_46, sout11_47, sout11_48,
    sout11_49, sout11_50, sout11_51, sout11_52, sout11_53, sout11_54, sout11_55, sout11_56, 
    sout11_57, sout11_58, sout11_59, sout11_60, sout11_61, sout11_62, sout11_63, sout11_64,
    
    sout12_1, sout12_2, sout12_3, sout12_4, sout12_5, sout12_6, sout12_7, sout12_8,
    sout12_9, sout12_10, sout12_11, sout12_12, sout12_13, sout12_14, sout12_15, sout12_16,
    sout12_17, sout12_18, sout12_19, sout12_20, sout12_21, sout12_22, sout12_23, sout12_24, 
    sout12_25, sout12_26, sout12_27, sout12_28, sout12_29, sout12_30, sout12_31, sout12_32,
    sout12_33, sout12_34, sout12_35, sout12_36, sout12_37, sout12_38, sout12_39, sout12_40,
    sout12_41, sout12_42, sout12_43, sout12_44, sout12_45, sout12_46, sout12_47, sout12_48,
    sout12_49, sout12_50, sout12_51, sout12_52, sout12_53, sout12_54, sout12_55, sout12_56, 
    sout12_57, sout12_58, sout12_59, sout12_60, sout12_61, sout12_62, sout12_63, sout12_64,
    
    sout13_1, sout13_2, sout13_3, sout13_4, sout13_5, sout13_6, sout13_7, sout13_8,
    sout13_9, sout13_10, sout13_11, sout13_12, sout13_13, sout13_14, sout13_15, sout13_16,
    sout13_17, sout13_18, sout13_19, sout13_20, sout13_21, sout13_22, sout13_23, sout13_24, 
    sout13_25, sout13_26, sout13_27, sout13_28, sout13_29, sout13_30, sout13_31, sout13_32,
    sout13_33, sout13_34, sout13_35, sout13_36, sout13_37, sout13_38, sout13_39, sout13_40,
    sout13_41, sout13_42, sout13_43, sout13_44, sout13_45, sout13_46, sout13_47, sout13_48,
    sout13_49, sout13_50, sout13_51, sout13_52, sout13_53, sout13_54, sout13_55, sout13_56, 
    sout13_57, sout13_58, sout13_59, sout13_60, sout13_61, sout13_62, sout13_63, sout13_64,
    
    sout14_1, sout14_2, sout14_3, sout14_4, sout14_5, sout14_6, sout14_7, sout14_8,
    sout14_9, sout14_10, sout14_11, sout14_12, sout14_13, sout14_14, sout14_15, sout14_16,
    sout14_17, sout14_18, sout14_19, sout14_20, sout14_21, sout14_22, sout14_23, sout14_24, 
    sout14_25, sout14_26, sout14_27, sout14_28, sout14_29, sout14_30, sout14_31, sout14_32,
    sout14_33, sout14_34, sout14_35, sout14_36, sout14_37, sout14_38, sout14_39, sout14_40,
    sout14_41, sout14_42, sout14_43, sout14_44, sout14_45, sout14_46, sout14_47, sout14_48,
    sout14_49, sout14_50, sout14_51, sout14_52, sout14_53, sout14_54, sout14_55, sout14_56, 
    sout14_57, sout14_58, sout14_59, sout14_60, sout14_61, sout14_62, sout14_63, sout14_64,
    
    sout15_1, sout15_2, sout15_3, sout15_4, sout15_5, sout15_6, sout15_7, sout15_8,
    sout15_9, sout15_10, sout15_11, sout15_12, sout15_13, sout15_14, sout15_15, sout15_16,
    sout15_17, sout15_18, sout15_19, sout15_20, sout15_21, sout15_22, sout15_23, sout15_24, 
    sout15_25, sout15_26, sout15_27, sout15_28, sout15_29, sout15_30, sout15_31, sout15_32,
    sout15_33, sout15_34, sout15_35, sout15_36, sout15_37, sout15_38, sout15_39, sout15_40,
    sout15_41, sout15_42, sout15_43, sout15_44, sout15_45, sout15_46, sout15_47, sout15_48,
    sout15_49, sout15_50, sout15_51, sout15_52, sout15_53, sout15_54, sout15_55, sout15_56, 
    sout15_57, sout15_58, sout15_59, sout15_60, sout15_61, sout15_62, sout15_63, sout15_64,
    
    sout16_1, sout16_2, sout16_3, sout16_4, sout16_5, sout16_6, sout16_7, sout16_8,
    sout16_9, sout16_10, sout16_11, sout16_12, sout16_13, sout16_14, sout16_15, sout16_16,
    sout16_17, sout16_18, sout16_19, sout16_20, sout16_21, sout16_22, sout16_23, sout16_24, 
    sout16_25, sout16_26, sout16_27, sout16_28, sout16_29, sout16_30, sout16_31, sout16_32,
    sout16_33, sout16_34, sout16_35, sout16_36, sout16_37, sout16_38, sout16_39, sout16_40,
    sout16_41, sout16_42, sout16_43, sout16_44, sout16_45, sout16_46, sout16_47, sout16_48,
    sout16_49, sout16_50, sout16_51, sout16_52, sout16_53, sout16_54, sout16_55, sout16_56, 
    sout16_57, sout16_58, sout16_59, sout16_60, sout16_61, sout16_62, sout16_63, sout16_64,
    
    sout17_1, sout17_2, sout17_3, sout17_4, sout17_5, sout17_6, sout17_7, sout17_8,
    sout17_9, sout17_10, sout17_11, sout17_12, sout17_13, sout17_14, sout17_15, sout17_16,
    sout17_17, sout17_18, sout17_19, sout17_20, sout17_21, sout17_22, sout17_23, sout17_24, 
    sout17_25, sout17_26, sout17_27, sout17_28, sout17_29, sout17_30, sout17_31, sout17_32,
    sout17_33, sout17_34, sout17_35, sout17_36, sout17_37, sout17_38, sout17_39, sout17_40,
    sout17_41, sout17_42, sout17_43, sout17_44, sout17_45, sout17_46, sout17_47, sout17_48,
    sout17_49, sout17_50, sout17_51, sout17_52, sout17_53, sout17_54, sout17_55, sout17_56, 
    sout17_57, sout17_58, sout17_59, sout17_60, sout17_61, sout17_62, sout17_63, sout17_64,
    
    sout18_1, sout18_2, sout18_3, sout18_4, sout18_5, sout18_6, sout18_7, sout18_8,
    sout18_9, sout18_10, sout18_11, sout18_12, sout18_13, sout18_14, sout18_15, sout18_16,
    sout18_17, sout18_18, sout18_19, sout18_20, sout18_21, sout18_22, sout18_23, sout18_24, 
    sout18_25, sout18_26, sout18_27, sout18_28, sout18_29, sout18_30, sout18_31, sout18_32,
    sout18_33, sout18_34, sout18_35, sout18_36, sout18_37, sout18_38, sout18_39, sout18_40,
    sout18_41, sout18_42, sout18_43, sout18_44, sout18_45, sout18_46, sout18_47, sout18_48,
    sout18_49, sout18_50, sout18_51, sout18_52, sout18_53, sout18_54, sout18_55, sout18_56, 
    sout18_57, sout18_58, sout18_59, sout18_60, sout18_61, sout18_62, sout18_63, sout18_64,
    
    sout19_1, sout19_2, sout19_3, sout19_4, sout19_5, sout19_6, sout19_7, sout19_8,
    sout19_9, sout19_10, sout19_11, sout19_12, sout19_13, sout19_14, sout19_15, sout19_16,
    sout19_17, sout19_18, sout19_19, sout19_20, sout19_21, sout19_22, sout19_23, sout19_24, 
    sout19_25, sout19_26, sout19_27, sout19_28, sout19_29, sout19_30, sout19_31, sout19_32,
    sout19_33, sout19_34, sout19_35, sout19_36, sout19_37, sout19_38, sout19_39, sout19_40,
    sout19_41, sout19_42, sout19_43, sout19_44, sout19_45, sout19_46, sout19_47, sout19_48,
    sout19_49, sout19_50, sout19_51, sout19_52, sout19_53, sout19_54, sout19_55, sout19_56, 
    sout19_57, sout19_58, sout19_59, sout19_60, sout19_61, sout19_62, sout19_63, sout19_64,
    
    sout20_1, sout20_2, sout20_3, sout20_4, sout20_5, sout20_6, sout20_7, sout20_8,
    sout20_9, sout20_10, sout20_11, sout20_12, sout20_13, sout20_14, sout20_15, sout20_16,
    sout20_17, sout20_18, sout20_19, sout20_20, sout20_21, sout20_22, sout20_23, sout20_24, 
    sout20_25, sout20_26, sout20_27, sout20_28, sout20_29, sout20_30, sout20_31, sout20_32,
    sout20_33, sout20_34, sout20_35, sout20_36, sout20_37, sout20_38, sout20_39, sout20_40,
    sout20_41, sout20_42, sout20_43, sout20_44, sout20_45, sout20_46, sout20_47, sout20_48,
    sout20_49, sout20_50, sout20_51, sout20_52, sout20_53, sout20_54, sout20_55, sout20_56, 
    sout20_57, sout20_58, sout20_59, sout20_60, sout20_61, sout20_62, sout20_63, sout20_64,
    
    sout21_1, sout21_2, sout21_3, sout21_4, sout21_5, sout21_6, sout21_7, sout21_8,
    sout21_9, sout21_10, sout21_11, sout21_12, sout21_13, sout21_14, sout21_15, sout21_16,
    sout21_17, sout21_18, sout21_19, sout21_20, sout21_21, sout21_22, sout21_23, sout21_24, 
    sout21_25, sout21_26, sout21_27, sout21_28, sout21_29, sout21_30, sout21_31, sout21_32,
    sout21_33, sout21_34, sout21_35, sout21_36, sout21_37, sout21_38, sout21_39, sout21_40,
    sout21_41, sout21_42, sout21_43, sout21_44, sout21_45, sout21_46, sout21_47, sout21_48,
    sout21_49, sout21_50, sout21_51, sout21_52, sout21_53, sout21_54, sout21_55, sout21_56, 
    sout21_57, sout21_58, sout21_59, sout21_60, sout21_61, sout21_62, sout21_63, sout21_64,
    
    sout22_1, sout22_2, sout22_3, sout22_4, sout22_5, sout22_6, sout22_7, sout22_8,
    sout22_9, sout22_10, sout22_11, sout22_12, sout22_13, sout22_14, sout22_15, sout22_16,
    sout22_17, sout22_18, sout22_19, sout22_20, sout22_21, sout22_22, sout22_23, sout22_24, 
    sout22_25, sout22_26, sout22_27, sout22_28, sout22_29, sout22_30, sout22_31, sout22_32,
    sout22_33, sout22_34, sout22_35, sout22_36, sout22_37, sout22_38, sout22_39, sout22_40,
    sout22_41, sout22_42, sout22_43, sout22_44, sout22_45, sout22_46, sout22_47, sout22_48,
    sout22_49, sout22_50, sout22_51, sout22_52, sout22_53, sout22_54, sout22_55, sout22_56, 
    sout22_57, sout22_58, sout22_59, sout22_60, sout22_61, sout22_62, sout22_63, sout22_64,
    
    sout23_1, sout23_2, sout23_3, sout23_4, sout23_5, sout23_6, sout23_7, sout23_8,
    sout23_9, sout23_10, sout23_11, sout23_12, sout23_13, sout23_14, sout23_15, sout23_16,
    sout23_17, sout23_18, sout23_19, sout23_20, sout23_21, sout23_22, sout23_23, sout23_24, 
    sout23_25, sout23_26, sout23_27, sout23_28, sout23_29, sout23_30, sout23_31, sout23_32,
    sout23_33, sout23_34, sout23_35, sout23_36, sout23_37, sout23_38, sout23_39, sout23_40,
    sout23_41, sout23_42, sout23_43, sout23_44, sout23_45, sout23_46, sout23_47, sout23_48,
    sout23_49, sout23_50, sout23_51, sout23_52, sout23_53, sout23_54, sout23_55, sout23_56, 
    sout23_57, sout23_58, sout23_59, sout23_60, sout23_61, sout23_62, sout23_63, sout23_64,
    
    sout24_1, sout24_2, sout24_3, sout24_4, sout24_5, sout24_6, sout24_7, sout24_8,
    sout24_9, sout24_10, sout24_11, sout24_12, sout24_13, sout24_14, sout24_15, sout24_16,
    sout24_17, sout24_18, sout24_19, sout24_20, sout24_21, sout24_22, sout24_23, sout24_24, 
    sout24_25, sout24_26, sout24_27, sout24_28, sout24_29, sout24_30, sout24_31, sout24_32,
    sout24_33, sout24_34, sout24_35, sout24_36, sout24_37, sout24_38, sout24_39, sout24_40,
    sout24_41, sout24_42, sout24_43, sout24_44, sout24_45, sout24_46, sout24_47, sout24_48,
    sout24_49, sout24_50, sout24_51, sout24_52, sout24_53, sout24_54, sout24_55, sout24_56, 
    sout24_57, sout24_58, sout24_59, sout24_60, sout24_61, sout24_62, sout24_63, sout24_64,
    
    sout25_1, sout25_2, sout25_3, sout25_4, sout25_5, sout25_6, sout25_7, sout25_8,
    sout25_9, sout25_10, sout25_11, sout25_12, sout25_13, sout25_14, sout25_15, sout25_16,
    sout25_17, sout25_18, sout25_19, sout25_20, sout25_21, sout25_22, sout25_23, sout25_24, 
    sout25_25, sout25_26, sout25_27, sout25_28, sout25_29, sout25_30, sout25_31, sout25_32,
    sout25_33, sout25_34, sout25_35, sout25_36, sout25_37, sout25_38, sout25_39, sout25_40,
    sout25_41, sout25_42, sout25_43, sout25_44, sout25_45, sout25_46, sout25_47, sout25_48,
    sout25_49, sout25_50, sout25_51, sout25_52, sout25_53, sout25_54, sout25_55, sout25_56, 
    sout25_57, sout25_58, sout25_59, sout25_60, sout25_61, sout25_62, sout25_63, sout25_64,
    
    sout26_1, sout26_2, sout26_3, sout26_4, sout26_5, sout26_6, sout26_7, sout26_8,
    sout26_9, sout26_10, sout26_11, sout26_12, sout26_13, sout26_14, sout26_15, sout26_16,
    sout26_17, sout26_18, sout26_19, sout26_20, sout26_21, sout26_22, sout26_23, sout26_24, 
    sout26_25, sout26_26, sout26_27, sout26_28, sout26_29, sout26_30, sout26_31, sout26_32,
    sout26_33, sout26_34, sout26_35, sout26_36, sout26_37, sout26_38, sout26_39, sout26_40,
    sout26_41, sout26_42, sout26_43, sout26_44, sout26_45, sout26_46, sout26_47, sout26_48,
    sout26_49, sout26_50, sout26_51, sout26_52, sout26_53, sout26_54, sout26_55, sout26_56, 
    sout26_57, sout26_58, sout26_59, sout26_60, sout26_61, sout26_62, sout26_63, sout26_64, 
    
    sout27_1, sout27_2, sout27_3, sout27_4, sout27_5, sout27_6, sout27_7, sout27_8,
    sout27_9, sout27_10, sout27_11, sout27_12, sout27_13, sout27_14, sout27_15, sout27_16,
    sout27_17, sout27_18, sout27_19, sout27_20, sout27_21, sout27_22, sout27_23, sout27_24, 
    sout27_25, sout27_26, sout27_27, sout27_28, sout27_29, sout27_30, sout27_31, sout27_32,
    sout27_33, sout27_34, sout27_35, sout27_36, sout27_37, sout27_38, sout27_39, sout27_40,
    sout27_41, sout27_42, sout27_43, sout27_44, sout27_45, sout27_46, sout27_47, sout27_48,
    sout27_49, sout27_50, sout27_51, sout27_52, sout27_53, sout27_54, sout27_55, sout27_56, 
    sout27_57, sout27_58, sout27_59, sout27_60, sout27_61, sout27_62, sout27_63, sout27_64,
    
    sout28_1, sout28_2, sout28_3, sout28_4, sout28_5, sout28_6, sout28_7, sout28_8,
    sout28_9, sout28_10, sout28_11, sout28_12, sout28_13, sout28_14, sout28_15, sout28_16,
    sout28_17, sout28_18, sout28_19, sout28_20, sout28_21, sout28_22, sout28_23, sout28_24, 
    sout28_25, sout28_26, sout28_27, sout28_28, sout28_29, sout28_30, sout28_31, sout28_32,
    sout28_33, sout28_34, sout28_35, sout28_36, sout28_37, sout28_38, sout28_39, sout28_40,
    sout28_41, sout28_42, sout28_43, sout28_44, sout28_45, sout28_46, sout28_47, sout28_48,
    sout28_49, sout28_50, sout28_51, sout28_52, sout28_53, sout28_54, sout28_55, sout28_56, 
    sout28_57, sout28_58, sout28_59, sout28_60, sout28_61, sout28_62, sout28_63, sout28_64,
    
    sout29_1, sout29_2, sout29_3, sout29_4, sout29_5, sout29_6, sout29_7, sout29_8,
    sout29_9, sout29_10, sout29_11, sout29_12, sout29_13, sout29_14, sout29_15, sout29_16,
    sout29_17, sout29_18, sout29_19, sout29_20, sout29_21, sout29_22, sout29_23, sout29_24, 
    sout29_25, sout29_26, sout29_27, sout29_28, sout29_29, sout29_30, sout29_31, sout29_32,
    sout29_33, sout29_34, sout29_35, sout29_36, sout29_37, sout29_38, sout29_39, sout29_40,
    sout29_41, sout29_42, sout29_43, sout29_44, sout29_45, sout29_46, sout29_47, sout29_48,
    sout29_49, sout29_50, sout29_51, sout29_52, sout29_53, sout29_54, sout29_55, sout29_56, 
    sout29_57, sout29_58, sout29_59, sout29_60, sout29_61, sout29_62, sout29_63, sout29_64,
    
    sout30_1, sout30_2, sout30_3, sout30_4, sout30_5, sout30_6, sout30_7, sout30_8,
    sout30_9, sout30_10, sout30_11, sout30_12, sout30_13, sout30_14, sout30_15, sout30_16,
    sout30_17, sout30_18, sout30_19, sout30_20, sout30_21, sout30_22, sout30_23, sout30_24, 
    sout30_25, sout30_26, sout30_27, sout30_28, sout30_29, sout30_30, sout30_31, sout30_32,
    sout30_33, sout30_34, sout30_35, sout30_36, sout30_37, sout30_38, sout30_39, sout30_40,
    sout30_41, sout30_42, sout30_43, sout30_44, sout30_45, sout30_46, sout30_47, sout30_48,
    sout30_49, sout30_50, sout30_51, sout30_52, sout30_53, sout30_54, sout30_55, sout30_56, 
    sout30_57, sout30_58, sout30_59, sout30_60, sout30_61, sout30_62, sout30_63, sout30_64,
    
    sout31_1, sout31_2, sout31_3, sout31_4, sout31_5, sout31_6, sout31_7, sout31_8,
    sout31_9, sout31_10, sout31_11, sout31_12, sout31_13, sout31_14, sout31_15, sout31_16,
    sout31_17, sout31_18, sout31_19, sout31_20, sout31_21, sout31_22, sout31_23, sout31_24, 
    sout31_25, sout31_26, sout31_27, sout31_28, sout31_29, sout31_30, sout31_31, sout31_32,
    sout31_33, sout31_34, sout31_35, sout31_36, sout31_37, sout31_38, sout31_39, sout31_40,
    sout31_41, sout31_42, sout31_43, sout31_44, sout31_45, sout31_46, sout31_47, sout31_48,
    sout31_49, sout31_50, sout31_51, sout31_52, sout31_53, sout31_54, sout31_55, sout31_56, 
    sout31_57, sout31_58, sout31_59, sout31_60, sout31_61, sout31_62, sout31_63, sout31_64,
    
    sout32_1, sout32_2, sout32_3, sout32_4, sout32_5, sout32_6, sout32_7, sout32_8,
    sout32_9, sout32_10, sout32_11, sout32_12, sout32_13, sout32_14, sout32_15, sout32_16,
    sout32_17, sout32_18, sout32_19, sout32_20, sout32_21, sout32_22, sout32_23, sout32_24, 
    sout32_25, sout32_26, sout32_27, sout32_28, sout32_29, sout32_30, sout32_31, sout32_32,
    sout32_33, sout32_34, sout32_35, sout32_36, sout32_37, sout32_38, sout32_39, sout32_40,
    sout32_41, sout32_42, sout32_43, sout32_44, sout32_45, sout32_46, sout32_47, sout32_48,
    sout32_49, sout32_50, sout32_51, sout32_52, sout32_53, sout32_54, sout32_55, sout32_56, 
    sout32_57, sout32_58, sout32_59, sout32_60, sout32_61, sout32_62, sout32_63, sout32_64,
    
    sout33_1, sout33_2, sout33_3, sout33_4, sout33_5, sout33_6, sout33_7, sout33_8,
    sout33_9, sout33_10, sout33_11, sout33_12, sout33_13, sout33_14, sout33_15, sout33_16,
    sout33_17, sout33_18, sout33_19, sout33_20, sout33_21, sout33_22, sout33_23, sout33_24, 
    sout33_25, sout33_26, sout33_27, sout33_28, sout33_29, sout33_30, sout33_31, sout33_32,
    sout33_33, sout33_34, sout33_35, sout33_36, sout33_37, sout33_38, sout33_39, sout33_40,
    sout33_41, sout33_42, sout33_43, sout33_44, sout33_45, sout33_46, sout33_47, sout33_48,
    sout33_49, sout33_50, sout33_51, sout33_52, sout33_53, sout33_54, sout33_55, sout33_56, 
    sout33_57, sout33_58, sout33_59, sout33_60, sout33_61, sout33_62, sout33_63, sout33_64,
                    
    sout34_1, sout34_2, sout34_3, sout34_4, sout34_5, sout34_6, sout34_7, sout34_8,
    sout34_9, sout34_10, sout34_11, sout34_12, sout34_13, sout34_14, sout34_15, sout34_16,
    sout34_17, sout34_18, sout34_19, sout34_20, sout34_21, sout34_22, sout34_23, sout34_24, 
    sout34_25, sout34_26, sout34_27, sout34_28, sout34_29, sout34_30, sout34_31, sout34_32,
    sout34_33, sout34_34, sout34_35, sout34_36, sout34_37, sout34_38, sout34_39, sout34_40,
    sout34_41, sout34_42, sout34_43, sout34_44, sout34_45, sout34_46, sout34_47, sout34_48,
    sout34_49, sout34_50, sout34_51, sout34_52, sout34_53, sout34_54, sout34_55, sout34_56, 
    sout34_57, sout34_58, sout34_59, sout34_60, sout34_61, sout34_62, sout34_63, sout34_64,
                  
    sout35_1, sout35_2, sout35_3, sout35_4, sout35_5, sout35_6, sout35_7, sout35_8,
    sout35_9, sout35_10, sout35_11, sout35_12, sout35_13, sout35_14, sout35_15, sout35_16,
    sout35_17, sout35_18, sout35_19, sout35_20, sout35_21, sout35_22, sout35_23, sout35_24, 
    sout35_25, sout35_26, sout35_27, sout35_28, sout35_29, sout35_30, sout35_31, sout35_32,
    sout35_33, sout35_34, sout35_35, sout35_36, sout35_37, sout35_38, sout35_39, sout35_40,
    sout35_41, sout35_42, sout35_43, sout35_44, sout35_45, sout35_46, sout35_47, sout35_48,
    sout35_49, sout35_50, sout35_51, sout35_52, sout35_53, sout35_54, sout35_55, sout35_56, 
    sout35_57, sout35_58, sout35_59, sout35_60, sout35_61, sout35_62, sout35_63, sout35_64,
                  
    sout36_1, sout36_2, sout36_3, sout36_4, sout36_5, sout36_6, sout36_7, sout36_8,
    sout36_9, sout36_10, sout36_11, sout36_12, sout36_13, sout36_14, sout36_15, sout36_16,
    sout36_17, sout36_18, sout36_19, sout36_20, sout36_21, sout36_22, sout36_23, sout36_24, 
    sout36_25, sout36_26, sout36_27, sout36_28, sout36_29, sout36_30, sout36_31, sout36_32,
    sout36_33, sout36_34, sout36_35, sout36_36, sout36_37, sout36_38, sout36_39, sout36_40,
    sout36_41, sout36_42, sout36_43, sout36_44, sout36_45, sout36_46, sout36_47, sout36_48,
    sout36_49, sout36_50, sout36_51, sout36_52, sout36_53, sout36_54, sout36_55, sout36_56, 
    sout36_57, sout36_58, sout36_59, sout36_60, sout36_61, sout36_62, sout36_63, sout36_64,
                  
    sout37_1, sout37_2, sout37_3, sout37_4, sout37_5, sout37_6, sout37_7, sout37_8,
    sout37_9, sout37_10, sout37_11, sout37_12, sout37_13, sout37_14, sout37_15, sout37_16,
    sout37_17, sout37_18, sout37_19, sout37_20, sout37_21, sout37_22, sout37_23, sout37_24, 
    sout37_25, sout37_26, sout37_27, sout37_28, sout37_29, sout37_30, sout37_31, sout37_32,
    sout37_33, sout37_34, sout37_35, sout37_36, sout37_37, sout37_38, sout37_39, sout37_40,
    sout37_41, sout37_42, sout37_43, sout37_44, sout37_45, sout37_46, sout37_47, sout37_48,
    sout37_49, sout37_50, sout37_51, sout37_52, sout37_53, sout37_54, sout37_55, sout37_56, 
    sout37_57, sout37_58, sout37_59, sout37_60, sout37_61, sout37_62, sout37_63, sout37_64,
                  
    sout38_1, sout38_2, sout38_3, sout38_4, sout38_5, sout38_6, sout38_7, sout38_8,
    sout38_9, sout38_10, sout38_11, sout38_12, sout38_13, sout38_14, sout38_15, sout38_16,
    sout38_17, sout38_18, sout38_19, sout38_20, sout38_21, sout38_22, sout38_23, sout38_24, 
    sout38_25, sout38_26, sout38_27, sout38_28, sout38_29, sout38_30, sout38_31, sout38_32,
    sout38_33, sout38_34, sout38_35, sout38_36, sout38_37, sout38_38, sout38_39, sout38_40,
    sout38_41, sout38_42, sout38_43, sout38_44, sout38_45, sout38_46, sout38_47, sout38_48,
    sout38_49, sout38_50, sout38_51, sout38_52, sout38_53, sout38_54, sout38_55, sout38_56, 
    sout38_57, sout38_58, sout38_59, sout38_60, sout38_61, sout38_62, sout38_63, sout38_64,
                  
    sout39_1, sout39_2, sout39_3, sout39_4, sout39_5, sout39_6, sout39_7, sout39_8,
    sout39_9, sout39_10, sout39_11, sout39_12, sout39_13, sout39_14, sout39_15, sout39_16,
    sout39_17, sout39_18, sout39_19, sout39_20, sout39_21, sout39_22, sout39_23, sout39_24, 
    sout39_25, sout39_26, sout39_27, sout39_28, sout39_29, sout39_30, sout39_31, sout39_32,
    sout39_33, sout39_34, sout39_35, sout39_36, sout39_37, sout39_38, sout39_39, sout39_40,
    sout39_41, sout39_42, sout39_43, sout39_44, sout39_45, sout39_46, sout39_47, sout39_48,
    sout39_49, sout39_50, sout39_51, sout39_52, sout39_53, sout39_54, sout39_55, sout39_56, 
    sout39_57, sout39_58, sout39_59, sout39_60, sout39_61, sout39_62, sout39_63, sout39_64,
                  
    sout40_1, sout40_2, sout40_3, sout40_4, sout40_5, sout40_6, sout40_7, sout40_8,
    sout40_9, sout40_10, sout40_11, sout40_12, sout40_13, sout40_14, sout40_15, sout40_16,
    sout40_17, sout40_18, sout40_19, sout40_20, sout40_21, sout40_22, sout40_23, sout40_24, 
    sout40_25, sout40_26, sout40_27, sout40_28, sout40_29, sout40_30, sout40_31, sout40_32,
    sout40_33, sout40_34, sout40_35, sout40_36, sout40_37, sout40_38, sout40_39, sout40_40,
    sout40_41, sout40_42, sout40_43, sout40_44, sout40_45, sout40_46, sout40_47, sout40_48,
    sout40_49, sout40_50, sout40_51, sout40_52, sout40_53, sout40_54, sout40_55, sout40_56, 
    sout40_57, sout40_58, sout40_59, sout40_60, sout40_61, sout40_62, sout40_63, sout40_64,
    
    sout41_1, sout41_2, sout41_3, sout41_4, sout41_5, sout41_6, sout41_7, sout41_8,
    sout41_9, sout41_10, sout41_11, sout41_12, sout41_13, sout41_14, sout41_15, sout41_16,
    sout41_17, sout41_18, sout41_19, sout41_20, sout41_21, sout41_22, sout41_23, sout41_24, 
    sout41_25, sout41_26, sout41_27, sout41_28, sout41_29, sout41_30, sout41_31, sout41_32,
    sout41_33, sout41_34, sout41_35, sout41_36, sout41_37, sout41_38, sout41_39, sout41_40,
    sout41_41, sout41_42, sout41_43, sout41_44, sout41_45, sout41_46, sout41_47, sout41_48,
    sout41_49, sout41_50, sout41_51, sout41_52, sout41_53, sout41_54, sout41_55, sout41_56, 
    sout41_57, sout41_58, sout41_59, sout41_60, sout41_61, sout41_62, sout41_63, sout41_64,
                  
    sout42_1, sout42_2, sout42_3, sout42_4, sout42_5, sout42_6, sout42_7, sout42_8,
    sout42_9, sout42_10, sout42_11, sout42_12, sout42_13, sout42_14, sout42_15, sout42_16,
    sout42_17, sout42_18, sout42_19, sout42_20, sout42_21, sout42_22, sout42_23, sout42_24, 
    sout42_25, sout42_26, sout42_27, sout42_28, sout42_29, sout42_30, sout42_31, sout42_32,
    sout42_33, sout42_34, sout42_35, sout42_36, sout42_37, sout42_38, sout42_39, sout42_40,
    sout42_41, sout42_42, sout42_43, sout42_44, sout42_45, sout42_46, sout42_47, sout42_48,
    sout42_49, sout42_50, sout42_51, sout42_52, sout42_53, sout42_54, sout42_55, sout42_56, 
    sout42_57, sout42_58, sout42_59, sout42_60, sout42_61, sout42_62, sout42_63, sout42_64,
                        
    sout43_1, sout43_2, sout43_3, sout43_4, sout43_5, sout43_6, sout43_7, sout43_8,
    sout43_9, sout43_10, sout43_11, sout43_12, sout43_13, sout43_14, sout43_15, sout43_16,
    sout43_17, sout43_18, sout43_19, sout43_20, sout43_21, sout43_22, sout43_23, sout43_24, 
    sout43_25, sout43_26, sout43_27, sout43_28, sout43_29, sout43_30, sout43_31, sout43_32,
    sout43_33, sout43_34, sout43_35, sout43_36, sout43_37, sout43_38, sout43_39, sout43_40,
    sout43_41, sout43_42, sout43_43, sout43_44, sout43_45, sout43_46, sout43_47, sout43_48,
    sout43_49, sout43_50, sout43_51, sout43_52, sout43_53, sout43_54, sout43_55, sout43_56, 
    sout43_57, sout43_58, sout43_59, sout43_60, sout43_61, sout43_62, sout43_63, sout43_64,
                  
    sout44_1, sout44_2, sout44_3, sout44_4, sout44_5, sout44_6, sout44_7, sout44_8,
    sout44_9, sout44_10, sout44_11, sout44_12, sout44_13, sout44_14, sout44_15, sout44_16,
    sout44_17, sout44_18, sout44_19, sout44_20, sout44_21, sout44_22, sout44_23, sout44_24, 
    sout44_25, sout44_26, sout44_27, sout44_28, sout44_29, sout44_30, sout44_31, sout44_32,
    sout44_33, sout44_34, sout44_35, sout44_36, sout44_37, sout44_38, sout44_39, sout44_40,
    sout44_41, sout44_42, sout44_43, sout44_44, sout44_45, sout44_46, sout44_47, sout44_48,
    sout44_49, sout44_50, sout44_51, sout44_52, sout44_53, sout44_54, sout44_55, sout44_56, 
    sout44_57, sout44_58, sout44_59, sout44_60, sout44_61, sout44_62, sout44_63, sout44_64,
                  
    sout45_1, sout45_2, sout45_3, sout45_4, sout45_5, sout45_6, sout45_7, sout45_8,
    sout45_9, sout45_10, sout45_11, sout45_12, sout45_13, sout45_14, sout45_15, sout45_16,
    sout45_17, sout45_18, sout45_19, sout45_20, sout45_21, sout45_22, sout45_23, sout45_24, 
    sout45_25, sout45_26, sout45_27, sout45_28, sout45_29, sout45_30, sout45_31, sout45_32,
    sout45_33, sout45_34, sout45_35, sout45_36, sout45_37, sout45_38, sout45_39, sout45_40,
    sout45_41, sout45_42, sout45_43, sout45_44, sout45_45, sout45_46, sout45_47, sout45_48,
    sout45_49, sout45_50, sout45_51, sout45_52, sout45_53, sout45_54, sout45_55, sout45_56, 
    sout45_57, sout45_58, sout45_59, sout45_60, sout45_61, sout45_62, sout45_63, sout45_64,
                  
    sout46_1, sout46_2, sout46_3, sout46_4, sout46_5, sout46_6, sout46_7, sout46_8,
    sout46_9, sout46_10, sout46_11, sout46_12, sout46_13, sout46_14, sout46_15, sout46_16,
    sout46_17, sout46_18, sout46_19, sout46_20, sout46_21, sout46_22, sout46_23, sout46_24, 
    sout46_25, sout46_26, sout46_27, sout46_28, sout46_29, sout46_30, sout46_31, sout46_32,
    sout46_33, sout46_34, sout46_35, sout46_36, sout46_37, sout46_38, sout46_39, sout46_40,
    sout46_41, sout46_42, sout46_43, sout46_44, sout46_45, sout46_46, sout46_47, sout46_48,
    sout46_49, sout46_50, sout46_51, sout46_52, sout46_53, sout46_54, sout46_55, sout46_56, 
    sout46_57, sout46_58, sout46_59, sout46_60, sout46_61, sout46_62, sout46_63, sout46_64,
                 
    sout47_1, sout47_2, sout47_3, sout47_4, sout47_5, sout47_6, sout47_7, sout47_8,
    sout47_9, sout47_10, sout47_11, sout47_12, sout47_13, sout47_14, sout47_15, sout47_16,
    sout47_17, sout47_18, sout47_19, sout47_20, sout47_21, sout47_22, sout47_23, sout47_24, 
    sout47_25, sout47_26, sout47_27, sout47_28, sout47_29, sout47_30, sout47_31, sout47_32,
    sout47_33, sout47_34, sout47_35, sout47_36, sout47_37, sout47_38, sout47_39, sout47_40,
    sout47_41, sout47_42, sout47_43, sout47_44, sout47_45, sout47_46, sout47_47, sout47_48,
    sout47_49, sout47_50, sout47_51, sout47_52, sout47_53, sout47_54, sout47_55, sout47_56, 
    sout47_57, sout47_58, sout47_59, sout47_60, sout47_61, sout47_62, sout47_63, sout47_64,
                  
    sout48_1, sout48_2, sout48_3, sout48_4, sout48_5, sout48_6, sout48_7, sout48_8,
    sout48_9, sout48_10, sout48_11, sout48_12, sout48_13, sout48_14, sout48_15, sout48_16,
    sout48_17, sout48_18, sout48_19, sout48_20, sout48_21, sout48_22, sout48_23, sout48_24, 
    sout48_25, sout48_26, sout48_27, sout48_28, sout48_29, sout48_30, sout48_31, sout48_32,
    sout48_33, sout48_34, sout48_35, sout48_36, sout48_37, sout48_38, sout48_39, sout48_40,
    sout48_41, sout48_42, sout48_43, sout48_44, sout48_45, sout48_46, sout48_47, sout48_48,
    sout48_49, sout48_50, sout48_51, sout48_52, sout48_53, sout48_54, sout48_55, sout48_56, 
    sout48_57, sout48_58, sout48_59, sout48_60, sout48_61, sout48_62, sout48_63, sout48_64,
                  
    sout49_1, sout49_2, sout49_3, sout49_4, sout49_5, sout49_6, sout49_7, sout49_8,
    sout49_9, sout49_10, sout49_11, sout49_12, sout49_13, sout49_14, sout49_15, sout49_16,
    sout49_17, sout49_18, sout49_19, sout49_20, sout49_21, sout49_22, sout49_23, sout49_24, 
    sout49_25, sout49_26, sout49_27, sout49_28, sout49_29, sout49_30, sout49_31, sout49_32,
    sout49_33, sout49_34, sout49_35, sout49_36, sout49_37, sout49_38, sout49_39, sout49_40,
    sout49_41, sout49_42, sout49_43, sout49_44, sout49_45, sout49_46, sout49_47, sout49_48,
    sout49_49, sout49_50, sout49_51, sout49_52, sout49_53, sout49_54, sout49_55, sout49_56, 
    sout49_57, sout49_58, sout49_59, sout49_60, sout49_61, sout49_62, sout49_63, sout49_64,
                  
    sout50_1, sout50_2, sout50_3, sout50_4, sout50_5, sout50_6, sout50_7, sout50_8,
    sout50_9, sout50_10, sout50_11, sout50_12, sout50_13, sout50_14, sout50_15, sout50_16,
    sout50_17, sout50_18, sout50_19, sout50_20, sout50_21, sout50_22, sout50_23, sout50_24, 
    sout50_25, sout50_26, sout50_27, sout50_28, sout50_29, sout50_30, sout50_31, sout50_32,
    sout50_33, sout50_34, sout50_35, sout50_36, sout50_37, sout50_38, sout50_39, sout50_40,
    sout50_41, sout50_42, sout50_43, sout50_44, sout50_45, sout50_46, sout50_47, sout50_48,
    sout50_49, sout50_50, sout50_51, sout50_52, sout50_53, sout50_54, sout50_55, sout50_56, 
    sout50_57, sout50_58, sout50_59, sout50_60, sout50_61, sout50_62, sout50_63, sout50_64,
    
    sout51_1, sout51_2, sout51_3, sout51_4, sout51_5, sout51_6, sout51_7, sout51_8,
    sout51_9, sout51_10, sout51_11, sout51_12, sout51_13, sout51_14, sout51_15, sout51_16,
    sout51_17, sout51_18, sout51_19, sout51_20, sout51_21, sout51_22, sout51_23, sout51_24, 
    sout51_25, sout51_26, sout51_27, sout51_28, sout51_29, sout51_30, sout51_31, sout51_32,
    sout51_33, sout51_34, sout51_35, sout51_36, sout51_37, sout51_38, sout51_39, sout51_40,
    sout51_41, sout51_42, sout51_43, sout51_44, sout51_45, sout51_46, sout51_47, sout51_48,
    sout51_49, sout51_50, sout51_51, sout51_52, sout51_53, sout51_54, sout51_55, sout51_56, 
    sout51_57, sout51_58, sout51_59, sout51_60, sout51_61, sout51_62, sout51_63, sout51_64,
                              
    sout52_1, sout52_2, sout52_3, sout52_4, sout52_5, sout52_6, sout52_7, sout52_8,
    sout52_9, sout52_10, sout52_11, sout52_12, sout52_13, sout52_14, sout52_15, sout52_16,
    sout52_17, sout52_18, sout52_19, sout52_20, sout52_21, sout52_22, sout52_23, sout52_24, 
    sout52_25, sout52_26, sout52_27, sout52_28, sout52_29, sout52_30, sout52_31, sout52_32,
    sout52_33, sout52_34, sout52_35, sout52_36, sout52_37, sout52_38, sout52_39, sout52_40,
    sout52_41, sout52_42, sout52_43, sout52_44, sout52_45, sout52_46, sout52_47, sout52_48,
    sout52_49, sout52_50, sout52_51, sout52_52, sout52_53, sout52_54, sout52_55, sout52_56, 
    sout52_57, sout52_58, sout52_59, sout52_60, sout52_61, sout52_62, sout52_63, sout52_64,
                  
    sout53_1, sout53_2, sout53_3, sout53_4, sout53_5, sout53_6, sout53_7, sout53_8,
    sout53_9, sout53_10, sout53_11, sout53_12, sout53_13, sout53_14, sout53_15, sout53_16,
    sout53_17, sout53_18, sout53_19, sout53_20, sout53_21, sout53_22, sout53_23, sout53_24, 
    sout53_25, sout53_26, sout53_27, sout53_28, sout53_29, sout53_30, sout53_31, sout53_32,
    sout53_33, sout53_34, sout53_35, sout53_36, sout53_37, sout53_38, sout53_39, sout53_40,
    sout53_41, sout53_42, sout53_43, sout53_44, sout53_45, sout53_46, sout53_47, sout53_48,
    sout53_49, sout53_50, sout53_51, sout53_52, sout53_53, sout53_54, sout53_55, sout53_56, 
    sout53_57, sout53_58, sout53_59, sout53_60, sout53_61, sout53_62, sout53_63, sout53_64,
                  
    sout54_1, sout54_2, sout54_3, sout54_4, sout54_5, sout54_6, sout54_7, sout54_8,
    sout54_9, sout54_10, sout54_11, sout54_12, sout54_13, sout54_14, sout54_15, sout54_16,
    sout54_17, sout54_18, sout54_19, sout54_20, sout54_21, sout54_22, sout54_23, sout54_24, 
    sout54_25, sout54_26, sout54_27, sout54_28, sout54_29, sout54_30, sout54_31, sout54_32,
    sout54_33, sout54_34, sout54_35, sout54_36, sout54_37, sout54_38, sout54_39, sout54_40,
    sout54_41, sout54_42, sout54_43, sout54_44, sout54_45, sout54_46, sout54_47, sout54_48,
    sout54_49, sout54_50, sout54_51, sout54_52, sout54_53, sout54_54, sout54_55, sout54_56, 
    sout54_57, sout54_58, sout54_59, sout54_60, sout54_61, sout54_62, sout54_63, sout54_64,
                  
    sout55_1, sout55_2, sout55_3, sout55_4, sout55_5, sout55_6, sout55_7, sout55_8,
    sout55_9, sout55_10, sout55_11, sout55_12, sout55_13, sout55_14, sout55_15, sout55_16,
    sout55_17, sout55_18, sout55_19, sout55_20, sout55_21, sout55_22, sout55_23, sout55_24, 
    sout55_25, sout55_26, sout55_27, sout55_28, sout55_29, sout55_30, sout55_31, sout55_32,
    sout55_33, sout55_34, sout55_35, sout55_36, sout55_37, sout55_38, sout55_39, sout55_40,
    sout55_41, sout55_42, sout55_43, sout55_44, sout55_45, sout55_46, sout55_47, sout55_48,
    sout55_49, sout55_50, sout55_51, sout55_52, sout55_53, sout55_54, sout55_55, sout55_56, 
    sout55_57, sout55_58, sout55_59, sout55_60, sout55_61, sout55_62, sout55_63, sout55_64,
                  
    sout56_1, sout56_2, sout56_3, sout56_4, sout56_5, sout56_6, sout56_7, sout56_8,
    sout56_9, sout56_10, sout56_11, sout56_12, sout56_13, sout56_14, sout56_15, sout56_16,
    sout56_17, sout56_18, sout56_19, sout56_20, sout56_21, sout56_22, sout56_23, sout56_24, 
    sout56_25, sout56_26, sout56_27, sout56_28, sout56_29, sout56_30, sout56_31, sout56_32,
    sout56_33, sout56_34, sout56_35, sout56_36, sout56_37, sout56_38, sout56_39, sout56_40,
    sout56_41, sout56_42, sout56_43, sout56_44, sout56_45, sout56_46, sout56_47, sout56_48,
    sout56_49, sout56_50, sout56_51, sout56_52, sout56_53, sout56_54, sout56_55, sout56_56, 
    sout56_57, sout56_58, sout56_59, sout56_60, sout56_61, sout56_62, sout56_63, sout56_64,
                  
    sout57_1, sout57_2, sout57_3, sout57_4, sout57_5, sout57_6, sout57_7, sout57_8,
    sout57_9, sout57_10, sout57_11, sout57_12, sout57_13, sout57_14, sout57_15, sout57_16,
    sout57_17, sout57_18, sout57_19, sout57_20, sout57_21, sout57_22, sout57_23, sout57_24, 
    sout57_25, sout57_26, sout57_27, sout57_28, sout57_29, sout57_30, sout57_31, sout57_32,
    sout57_33, sout57_34, sout57_35, sout57_36, sout57_37, sout57_38, sout57_39, sout57_40,
    sout57_41, sout57_42, sout57_43, sout57_44, sout57_45, sout57_46, sout57_47, sout57_48,
    sout57_49, sout57_50, sout57_51, sout57_52, sout57_53, sout57_54, sout57_55, sout57_56, 
    sout57_57, sout57_58, sout57_59, sout57_60, sout57_61, sout57_62, sout57_63, sout57_64,
                  
    sout58_1, sout58_2, sout58_3, sout58_4, sout58_5, sout58_6, sout58_7, sout58_8,
    sout58_9, sout58_10, sout58_11, sout58_12, sout58_13, sout58_14, sout58_15, sout58_16,
    sout58_17, sout58_18, sout58_19, sout58_20, sout58_21, sout58_22, sout58_23, sout58_24, 
    sout58_25, sout58_26, sout58_27, sout58_28, sout58_29, sout58_30, sout58_31, sout58_32,
    sout58_33, sout58_34, sout58_35, sout58_36, sout58_37, sout58_38, sout58_39, sout58_40,
    sout58_41, sout58_42, sout58_43, sout58_44, sout58_45, sout58_46, sout58_47, sout58_48,
    sout58_49, sout58_50, sout58_51, sout58_52, sout58_53, sout58_54, sout58_55, sout58_56, 
    sout58_57, sout58_58, sout58_59, sout58_60, sout58_61, sout58_62, sout58_63, sout58_64,
                  
    sout59_1, sout59_2, sout59_3, sout59_4, sout59_5, sout59_6, sout59_7, sout59_8,
    sout59_9, sout59_10, sout59_11, sout59_12, sout59_13, sout59_14, sout59_15, sout59_16,
    sout59_17, sout59_18, sout59_19, sout59_20, sout59_21, sout59_22, sout59_23, sout59_24, 
    sout59_25, sout59_26, sout59_27, sout59_28, sout59_29, sout59_30, sout59_31, sout59_32,
    sout59_33, sout59_34, sout59_35, sout59_36, sout59_37, sout59_38, sout59_39, sout59_40,
    sout59_41, sout59_42, sout59_43, sout59_44, sout59_45, sout59_46, sout59_47, sout59_48,
    sout59_49, sout59_50, sout59_51, sout59_52, sout59_53, sout59_54, sout59_55, sout59_56, 
    sout59_57, sout59_58, sout59_59, sout59_60, sout59_61, sout59_62, sout59_63, sout59_64,
                  
    sout60_1, sout60_2, sout60_3, sout60_4, sout60_5, sout60_6, sout60_7, sout60_8,
    sout60_9, sout60_10, sout60_11, sout60_12, sout60_13, sout60_14, sout60_15, sout60_16,
    sout60_17, sout60_18, sout60_19, sout60_20, sout60_21, sout60_22, sout60_23, sout60_24, 
    sout60_25, sout60_26, sout60_27, sout60_28, sout60_29, sout60_30, sout60_31, sout60_32,
    sout60_33, sout60_34, sout60_35, sout60_36, sout60_37, sout60_38, sout60_39, sout60_40,
    sout60_41, sout60_42, sout60_43, sout60_44, sout60_45, sout60_46, sout60_47, sout60_48,
    sout60_49, sout60_50, sout60_51, sout60_52, sout60_53, sout60_54, sout60_55, sout60_56, 
    sout60_57, sout60_58, sout60_59, sout60_60, sout60_61, sout60_62, sout60_63, sout60_64,
                  
    sout61_1, sout61_2, sout61_3, sout61_4, sout61_5, sout61_6, sout61_7, sout61_8,
    sout61_9, sout61_10, sout61_11, sout61_12, sout61_13, sout61_14, sout61_15, sout61_16,
    sout61_17, sout61_18, sout61_19, sout61_20, sout61_21, sout61_22, sout61_23, sout61_24, 
    sout61_25, sout61_26, sout61_27, sout61_28, sout61_29, sout61_30, sout61_31, sout61_32,
    sout61_33, sout61_34, sout61_35, sout61_36, sout61_37, sout61_38, sout61_39, sout61_40,
    sout61_41, sout61_42, sout61_43, sout61_44, sout61_45, sout61_46, sout61_47, sout61_48,
    sout61_49, sout61_50, sout61_51, sout61_52, sout61_53, sout61_54, sout61_55, sout61_56, 
    sout61_57, sout61_58, sout61_59, sout61_60, sout61_61, sout61_62, sout61_63, sout61_64,
                  
    sout62_1, sout62_2, sout62_3, sout62_4, sout62_5, sout62_6, sout62_7, sout62_8,
    sout62_9, sout62_10, sout62_11, sout62_12, sout62_13, sout62_14, sout62_15, sout62_16,
    sout62_17, sout62_18, sout62_19, sout62_20, sout62_21, sout62_22, sout62_23, sout62_24, 
    sout62_25, sout62_26, sout62_27, sout62_28, sout62_29, sout62_30, sout62_31, sout62_32,
    sout62_33, sout62_34, sout62_35, sout62_36, sout62_37, sout62_38, sout62_39, sout62_40,
    sout62_41, sout62_42, sout62_43, sout62_44, sout62_45, sout62_46, sout62_47, sout62_48,
    sout62_49, sout62_50, sout62_51, sout62_52, sout62_53, sout62_54, sout62_55, sout62_56, 
    sout62_57, sout62_58, sout62_59, sout62_60, sout62_61, sout62_62, sout62_63, sout62_64,
                  
    sout63_1, sout63_2, sout63_3, sout63_4, sout63_5, sout63_6, sout63_7, sout63_8,
    sout63_9, sout63_10, sout63_11, sout63_12, sout63_13, sout63_14, sout63_15, sout63_16,
    sout63_17, sout63_18, sout63_19, sout63_20, sout63_21, sout63_22, sout63_23, sout63_24, 
    sout63_25, sout63_26, sout63_27, sout63_28, sout63_29, sout63_30, sout63_31, sout63_32,
    sout63_33, sout63_34, sout63_35, sout63_36, sout63_37, sout63_38, sout63_39, sout63_40,
    sout63_41, sout63_42, sout63_43, sout63_44, sout63_45, sout63_46, sout63_47, sout63_48,
    sout63_49, sout63_50, sout63_51, sout63_52, sout63_53, sout63_54, sout63_55, sout63_56, 
    sout63_57, sout63_58, sout63_59, sout63_60, sout63_61, sout63_62, sout63_63, sout63_64,
                  
    sout64_1, sout64_2, sout64_3, sout64_4, sout64_5, sout64_6, sout64_7, sout64_8,
    sout64_9, sout64_10, sout64_11, sout64_12, sout64_13, sout64_14, sout64_15, sout64_16,
    sout64_17, sout64_18, sout64_19, sout64_20, sout64_21, sout64_22, sout64_23, sout64_24, 
    sout64_25, sout64_26, sout64_27, sout64_28, sout64_29, sout64_30, sout64_31, sout64_32,
    sout64_33, sout64_34, sout64_35, sout64_36, sout64_37, sout64_38, sout64_39, sout64_40,
    sout64_41, sout64_42, sout64_43, sout64_44, sout64_45, sout64_46, sout64_47, sout64_48,
    sout64_49, sout64_50, sout64_51, sout64_52, sout64_53, sout64_54, sout64_55, sout64_56, 
    sout64_57, sout64_58, sout64_59, sout64_60, sout64_61, sout64_62, sout64_63, sout64_64    
    );
    
    input clk, rst;
    
    input [7:0] ain1, ain2, ain3, ain4, ain5, ain6, ain7, ain8,
                ain9, ain10, ain11, ain12, ain13, ain14, ain15, ain16, 
                ain17, ain18, ain19, ain20, ain21, ain22, ain23, ain24, 
                ain25, ain26, ain27, ain28, ain29, ain30, ain31, ain32, 
                ain33, ain34, ain35, ain36, ain37, ain38, ain39, ain40, 
                ain41, ain42, ain43, ain44, ain45, ain46, ain47, ain48,
                ain49, ain50, ain51, ain52, ain53, ain54, ain55, ain56,
                ain57, ain58, ain59, ain60, ain61, ain62, ain63, ain64;
                
    input [7:0] win1, win2, win3, win4, win5, win6, win7, win8,
                win9, win10, win11, win12, win13, win14, win15, win16, 
                win17, win18, win19, win20, win21, win22, win23, win24, 
                win25, win26, win27, win28, win29, win30, win31, win32, 
                win33, win34, win35, win36, win37, win38, win39, win40, 
                win41, win42, win43, win44, win45, win46, win47, win48,
                win49, win50, win51, win52, win53, win54, win55, win56,
                win57, win58, win59, win60, win61, win62, win63, win64;  
                
    //row1
    output [21:0] sout11, sout12, sout13, sout14, sout15, sout16, sout17, sout18,
                  sout19, sout1_10, sout1_11, sout1_12, sout1_13, sout1_14, sout1_15, sout1_16,
                  sout1_17, sout1_18, sout1_19, sout1_20, sout1_21, sout1_22, sout1_23, sout1_24, 
                  sout1_25, sout1_26, sout1_27, sout1_28, sout1_29, sout1_30, sout1_31, sout1_32,
                  sout1_33, sout1_34, sout1_35, sout1_36, sout1_37, sout1_38, sout1_39, sout1_40,
                  sout1_41, sout1_42, sout1_43, sout1_44, sout1_45, sout1_46, sout1_47, sout1_48,
                  sout1_49, sout1_50, sout1_51, sout1_52, sout1_53, sout1_54, sout1_55, sout1_56, 
                  sout1_57, sout1_58, sout1_59, sout1_60, sout1_61, sout1_62, sout1_63, sout1_64;
    
    //row2       
    output [21:0] sout21, sout22, sout23, sout24, sout25, sout26, sout27, sout28,
                  sout29, sout2_10, sout2_11, sout2_12, sout2_13, sout2_14, sout2_15, sout2_16,
                  sout2_17, sout2_18, sout2_19, sout2_20, sout2_21, sout2_22, sout2_23, sout2_24, 
                  sout2_25, sout2_26, sout2_27, sout2_28, sout2_29, sout2_30, sout2_31, sout2_32,
                  sout2_33, sout2_34, sout2_35, sout2_36, sout2_37, sout2_38, sout2_39, sout2_40,
                  sout2_41, sout2_42, sout2_43, sout2_44, sout2_45, sout2_46, sout2_47, sout2_48,
                  sout2_49, sout2_50, sout2_51, sout2_52, sout2_53, sout2_54, sout2_55, sout2_56, 
                  sout2_57, sout2_58, sout2_59, sout2_60, sout2_61, sout2_62, sout2_63, sout2_64;
        
    //row3          
    output [21:0] sout31, sout32, sout33, sout34, sout35, sout36, sout37, sout38,
                  sout39, sout3_10, sout3_11, sout3_12, sout3_13, sout3_14, sout3_15, sout3_16,
                  sout3_17, sout3_18, sout3_19, sout3_20, sout3_21, sout3_22, sout3_23, sout3_24, 
                  sout3_25, sout3_26, sout3_27, sout3_28, sout3_29, sout3_30, sout3_31, sout3_32,
                  sout3_33, sout3_34, sout3_35, sout3_36, sout3_37, sout3_38, sout3_39, sout3_40,
                  sout3_41, sout3_42, sout3_43, sout3_44, sout3_45, sout3_46, sout3_47, sout3_48,
                  sout3_49, sout3_50, sout3_51, sout3_52, sout3_53, sout3_54, sout3_55, sout3_56, 
                  sout3_57, sout3_58, sout3_59, sout3_60, sout3_61, sout3_62, sout3_63, sout3_64;
                
    //row4                
    output [21:0] sout41, sout42, sout43, sout44, sout45, sout46, sout47, sout48,
                  sout49, sout4_10, sout4_11, sout4_12, sout4_13, sout4_14, sout4_15, sout4_16,
                  sout4_17, sout4_18, sout4_19, sout4_20, sout4_21, sout4_22, sout4_23, sout4_24, 
                  sout4_25, sout4_26, sout4_27, sout4_28, sout4_29, sout4_30, sout4_31, sout4_32,
                  sout4_33, sout4_34, sout4_35, sout4_36, sout4_37, sout4_38, sout4_39, sout4_40,
                  sout4_41, sout4_42, sout4_43, sout4_44, sout4_45, sout4_46, sout4_47, sout4_48,
                  sout4_49, sout4_50, sout4_51, sout4_52, sout4_53, sout4_54, sout4_55, sout4_56, 
                  sout4_57, sout4_58, sout4_59, sout4_60, sout4_61, sout4_62, sout4_63, sout4_64;
           
    //row5               
    output [21:0] sout51, sout52, sout53, sout54, sout55, sout56, sout57, sout58,
                  sout59, sout5_10, sout5_11, sout5_12, sout5_13, sout5_14, sout5_15, sout5_16,
                  sout5_17, sout5_18, sout5_19, sout5_20, sout5_21, sout5_22, sout5_23, sout5_24, 
                  sout5_25, sout5_26, sout5_27, sout5_28, sout5_29, sout5_30, sout5_31, sout5_32,
                  sout5_33, sout5_34, sout5_35, sout5_36, sout5_37, sout5_38, sout5_39, sout5_40,
                  sout5_41, sout5_42, sout5_43, sout5_44, sout5_45, sout5_46, sout5_47, sout5_48,
                  sout5_49, sout5_50, sout5_51, sout5_52, sout5_53, sout5_54, sout5_55, sout5_56, 
                  sout5_57, sout5_58, sout5_59, sout5_60, sout5_61, sout5_62, sout5_63, sout5_64;
         
    //row6         
    output [21:0] sout61, sout62, sout63, sout64, sout65, sout66, sout67, sout68,
                  sout69, sout6_10, sout6_11, sout6_12, sout6_13, sout6_14, sout6_15, sout6_16,
                  sout6_17, sout6_18, sout6_19, sout6_20, sout6_21, sout6_22, sout6_23, sout6_24, 
                  sout6_25, sout6_26, sout6_27, sout6_28, sout6_29, sout6_30, sout6_31, sout6_32,
                  sout6_33, sout6_34, sout6_35, sout6_36, sout6_37, sout6_38, sout6_39, sout6_40,
                  sout6_41, sout6_42, sout6_43, sout6_44, sout6_45, sout6_46, sout6_47, sout6_48,
                  sout6_49, sout6_50, sout6_51, sout6_52, sout6_53, sout6_54, sout6_55, sout6_56, 
                  sout6_57, sout6_58, sout6_59, sout6_60, sout6_61, sout6_62, sout6_63, sout6_64;
              
    //row7    
    output [21:0] sout71, sout72, sout73, sout74, sout75, sout76, sout77, sout78,
                  sout79, sout7_10, sout7_11, sout7_12, sout7_13, sout7_14, sout7_15, sout7_16,
                  sout7_17, sout7_18, sout7_19, sout7_20, sout7_21, sout7_22, sout7_23, sout7_24, 
                  sout7_25, sout7_26, sout7_27, sout7_28, sout7_29, sout7_30, sout7_31, sout7_32,
                  sout7_33, sout7_34, sout7_35, sout7_36, sout7_37, sout7_38, sout7_39, sout7_40,
                  sout7_41, sout7_42, sout7_43, sout7_44, sout7_45, sout7_46, sout7_47, sout7_48,
                  sout7_49, sout7_50, sout7_51, sout7_52, sout7_53, sout7_54, sout7_55, sout7_56, 
                  sout7_57, sout7_58, sout7_59, sout7_60, sout7_61, sout7_62, sout7_63, sout7_64;
              
    //row8    
    output [21:0] sout81, sout82, sout83, sout84, sout85, sout86, sout87, sout88,
                  sout89, sout8_10, sout8_11, sout8_12, sout8_13, sout8_14, sout8_15, sout8_16,
                  sout8_17, sout8_18, sout8_19, sout8_20, sout8_21, sout8_22, sout8_23, sout8_24, 
                  sout8_25, sout8_26, sout8_27, sout8_28, sout8_29, sout8_30, sout8_31, sout8_32,
                  sout8_33, sout8_34, sout8_35, sout8_36, sout8_37, sout8_38, sout8_39, sout8_40,
                  sout8_41, sout8_42, sout8_43, sout8_44, sout8_45, sout8_46, sout8_47, sout8_48,
                  sout8_49, sout8_50, sout8_51, sout8_52, sout8_53, sout8_54, sout8_55, sout8_56, 
                  sout8_57, sout8_58, sout8_59, sout8_60, sout8_61, sout8_62, sout8_63, sout8_64;
        
    //row9                
    output [21:0] sout91, sout92, sout93, sout94, sout95, sout96, sout97, sout98,
                  sout99, sout9_10, sout9_11, sout9_12, sout9_13, sout9_14, sout9_15, sout9_16,
                  sout9_17, sout9_18, sout9_19, sout9_20, sout9_21, sout9_22, sout9_23, sout9_24, 
                  sout9_25, sout9_26, sout9_27, sout9_28, sout9_29, sout9_30, sout9_31, sout9_32,
                  sout9_33, sout9_34, sout9_35, sout9_36, sout9_37, sout9_38, sout9_39, sout9_40,
                  sout9_41, sout9_42, sout9_43, sout9_44, sout9_45, sout9_46, sout9_47, sout9_48,
                  sout9_49, sout9_50, sout9_51, sout9_52, sout9_53, sout9_54, sout9_55, sout9_56, 
                  sout9_57, sout9_58, sout9_59, sout9_60, sout9_61, sout9_62, sout9_63, sout9_64;
           
    //row10 
    output [21:0] sout10_1, sout10_2, sout10_3, sout10_4, sout10_5, sout10_6, sout10_7, sout10_8,
                  sout10_9, sout10_10, sout10_11, sout10_12, sout10_13, sout10_14, sout10_15, sout10_16,
                  sout10_17, sout10_18, sout10_19, sout10_20, sout10_21, sout10_22, sout10_23, sout10_24, 
                  sout10_25, sout10_26, sout10_27, sout10_28, sout10_29, sout10_30, sout10_31, sout10_32,
                  sout10_33, sout10_34, sout10_35, sout10_36, sout10_37, sout10_38, sout10_39, sout10_40,
                  sout10_41, sout10_42, sout10_43, sout10_44, sout10_45, sout10_46, sout10_47, sout10_48,
                  sout10_49, sout10_50, sout10_51, sout10_52, sout10_53, sout10_54, sout10_55, sout10_56, 
                  sout10_57, sout10_58, sout10_59, sout10_60, sout10_61, sout10_62, sout10_63, sout10_64;
                  
    //row11
    output [21:0] sout11_1, sout11_2, sout11_3, sout11_4, sout11_5, sout11_6, sout11_7, sout11_8,
                  sout11_9, sout11_10, sout11_11, sout11_12, sout11_13, sout11_14, sout11_15, sout11_16,
                  sout11_17, sout11_18, sout11_19, sout11_20, sout11_21, sout11_22, sout11_23, sout11_24, 
                  sout11_25, sout11_26, sout11_27, sout11_28, sout11_29, sout11_30, sout11_31, sout11_32,
                  sout11_33, sout11_34, sout11_35, sout11_36, sout11_37, sout11_38, sout11_39, sout11_40,
                  sout11_41, sout11_42, sout11_43, sout11_44, sout11_45, sout11_46, sout11_47, sout11_48,
                  sout11_49, sout11_50, sout11_51, sout11_52, sout11_53, sout11_54, sout11_55, sout11_56, 
                  sout11_57, sout11_58, sout11_59, sout11_60, sout11_61, sout11_62, sout11_63, sout11_64;
                        
    //row12
    output [21:0] sout12_1, sout12_2, sout12_3, sout12_4, sout12_5, sout12_6, sout12_7, sout12_8,
                  sout12_9, sout12_10, sout12_11, sout12_12, sout12_13, sout12_14, sout12_15, sout12_16,
                  sout12_17, sout12_18, sout12_19, sout12_20, sout12_21, sout12_22, sout12_23, sout12_24, 
                  sout12_25, sout12_26, sout12_27, sout12_28, sout12_29, sout12_30, sout12_31, sout12_32,
                  sout12_33, sout12_34, sout12_35, sout12_36, sout12_37, sout12_38, sout12_39, sout12_40,
                  sout12_41, sout12_42, sout12_43, sout12_44, sout12_45, sout12_46, sout12_47, sout12_48,
                  sout12_49, sout12_50, sout12_51, sout12_52, sout12_53, sout12_54, sout12_55, sout12_56, 
                  sout12_57, sout12_58, sout12_59, sout12_60, sout12_61, sout12_62, sout12_63, sout12_64;
                  
    //row13
    output [21:0] sout13_1, sout13_2, sout13_3, sout13_4, sout13_5, sout13_6, sout13_7, sout13_8,
                  sout13_9, sout13_10, sout13_11, sout13_12, sout13_13, sout13_14, sout13_15, sout13_16,
                  sout13_17, sout13_18, sout13_19, sout13_20, sout13_21, sout13_22, sout13_23, sout13_24, 
                  sout13_25, sout13_26, sout13_27, sout13_28, sout13_29, sout13_30, sout13_31, sout13_32,
                  sout13_33, sout13_34, sout13_35, sout13_36, sout13_37, sout13_38, sout13_39, sout13_40,
                  sout13_41, sout13_42, sout13_43, sout13_44, sout13_45, sout13_46, sout13_47, sout13_48,
                  sout13_49, sout13_50, sout13_51, sout13_52, sout13_53, sout13_54, sout13_55, sout13_56, 
                  sout13_57, sout13_58, sout13_59, sout13_60, sout13_61, sout13_62, sout13_63, sout13_64;
                  
    //row14
    output [21:0] sout14_1, sout14_2, sout14_3, sout14_4, sout14_5, sout14_6, sout14_7, sout14_8,
                  sout14_9, sout14_10, sout14_11, sout14_12, sout14_13, sout14_14, sout14_15, sout14_16,
                  sout14_17, sout14_18, sout14_19, sout14_20, sout14_21, sout14_22, sout14_23, sout14_24, 
                  sout14_25, sout14_26, sout14_27, sout14_28, sout14_29, sout14_30, sout14_31, sout14_32,
                  sout14_33, sout14_34, sout14_35, sout14_36, sout14_37, sout14_38, sout14_39, sout14_40,
                  sout14_41, sout14_42, sout14_43, sout14_44, sout14_45, sout14_46, sout14_47, sout14_48,
                  sout14_49, sout14_50, sout14_51, sout14_52, sout14_53, sout14_54, sout14_55, sout14_56, 
                  sout14_57, sout14_58, sout14_59, sout14_60, sout14_61, sout14_62, sout14_63, sout14_64;
                  
    //row15
    output [21:0] sout15_1, sout15_2, sout15_3, sout15_4, sout15_5, sout15_6, sout15_7, sout15_8,
                  sout15_9, sout15_10, sout15_11, sout15_12, sout15_13, sout15_14, sout15_15, sout15_16,
                  sout15_17, sout15_18, sout15_19, sout15_20, sout15_21, sout15_22, sout15_23, sout15_24, 
                  sout15_25, sout15_26, sout15_27, sout15_28, sout15_29, sout15_30, sout15_31, sout15_32,
                  sout15_33, sout15_34, sout15_35, sout15_36, sout15_37, sout15_38, sout15_39, sout15_40,
                  sout15_41, sout15_42, sout15_43, sout15_44, sout15_45, sout15_46, sout15_47, sout15_48,
                  sout15_49, sout15_50, sout15_51, sout15_52, sout15_53, sout15_54, sout15_55, sout15_56, 
                  sout15_57, sout15_58, sout15_59, sout15_60, sout15_61, sout15_62, sout15_63, sout15_64;
                  
    //row16
    output [21:0] sout16_1, sout16_2, sout16_3, sout16_4, sout16_5, sout16_6, sout16_7, sout16_8,
                  sout16_9, sout16_10, sout16_11, sout16_12, sout16_13, sout16_14, sout16_15, sout16_16,
                  sout16_17, sout16_18, sout16_19, sout16_20, sout16_21, sout16_22, sout16_23, sout16_24, 
                  sout16_25, sout16_26, sout16_27, sout16_28, sout16_29, sout16_30, sout16_31, sout16_32,
                  sout16_33, sout16_34, sout16_35, sout16_36, sout16_37, sout16_38, sout16_39, sout16_40,
                  sout16_41, sout16_42, sout16_43, sout16_44, sout16_45, sout16_46, sout16_47, sout16_48,
                  sout16_49, sout16_50, sout16_51, sout16_52, sout16_53, sout16_54, sout16_55, sout16_56, 
                  sout16_57, sout16_58, sout16_59, sout16_60, sout16_61, sout16_62, sout16_63, sout16_64;
                
    //row17
    output [21:0] sout17_1, sout17_2, sout17_3, sout17_4, sout17_5, sout17_6, sout17_7, sout17_8,
                  sout17_9, sout17_10, sout17_11, sout17_12, sout17_13, sout17_14, sout17_15, sout17_16,
                  sout17_17, sout17_18, sout17_19, sout17_20, sout17_21, sout17_22, sout17_23, sout17_24, 
                  sout17_25, sout17_26, sout17_27, sout17_28, sout17_29, sout17_30, sout17_31, sout17_32,
                  sout17_33, sout17_34, sout17_35, sout17_36, sout17_37, sout17_38, sout17_39, sout17_40,
                  sout17_41, sout17_42, sout17_43, sout17_44, sout17_45, sout17_46, sout17_47, sout17_48,
                  sout17_49, sout17_50, sout17_51, sout17_52, sout17_53, sout17_54, sout17_55, sout17_56, 
                  sout17_57, sout17_58, sout17_59, sout17_60, sout17_61, sout17_62, sout17_63, sout17_64;
                  
    //row18
    output [21:0] sout18_1, sout18_2, sout18_3, sout18_4, sout18_5, sout18_6, sout18_7, sout18_8,
                  sout18_9, sout18_10, sout18_11, sout18_12, sout18_13, sout18_14, sout18_15, sout18_16,
                  sout18_17, sout18_18, sout18_19, sout18_20, sout18_21, sout18_22, sout18_23, sout18_24, 
                  sout18_25, sout18_26, sout18_27, sout18_28, sout18_29, sout18_30, sout18_31, sout18_32,
                  sout18_33, sout18_34, sout18_35, sout18_36, sout18_37, sout18_38, sout18_39, sout18_40,
                  sout18_41, sout18_42, sout18_43, sout18_44, sout18_45, sout18_46, sout18_47, sout18_48,
                  sout18_49, sout18_50, sout18_51, sout18_52, sout18_53, sout18_54, sout18_55, sout18_56, 
                  sout18_57, sout18_58, sout18_59, sout18_60, sout18_61, sout18_62, sout18_63, sout18_64;
                  
    //row19
    output [21:0] sout19_1, sout19_2, sout19_3, sout19_4, sout19_5, sout19_6, sout19_7, sout19_8,
                  sout19_9, sout19_10, sout19_11, sout19_12, sout19_13, sout19_14, sout19_15, sout19_16,
                  sout19_17, sout19_18, sout19_19, sout19_20, sout19_21, sout19_22, sout19_23, sout19_24, 
                  sout19_25, sout19_26, sout19_27, sout19_28, sout19_29, sout19_30, sout19_31, sout19_32,
                  sout19_33, sout19_34, sout19_35, sout19_36, sout19_37, sout19_38, sout19_39, sout19_40,
                  sout19_41, sout19_42, sout19_43, sout19_44, sout19_45, sout19_46, sout19_47, sout19_48,
                  sout19_49, sout19_50, sout19_51, sout19_52, sout19_53, sout19_54, sout19_55, sout19_56, 
                  sout19_57, sout19_58, sout19_59, sout19_60, sout19_61, sout19_62, sout19_63, sout19_64;
                  
    //row20
    output [21:0] sout20_1, sout20_2, sout20_3, sout20_4, sout20_5, sout20_6, sout20_7, sout20_8,
                  sout20_9, sout20_10, sout20_11, sout20_12, sout20_13, sout20_14, sout20_15, sout20_16,
                  sout20_17, sout20_18, sout20_19, sout20_20, sout20_21, sout20_22, sout20_23, sout20_24, 
                  sout20_25, sout20_26, sout20_27, sout20_28, sout20_29, sout20_30, sout20_31, sout20_32,
                  sout20_33, sout20_34, sout20_35, sout20_36, sout20_37, sout20_38, sout20_39, sout20_40,
                  sout20_41, sout20_42, sout20_43, sout20_44, sout20_45, sout20_46, sout20_47, sout20_48,
                  sout20_49, sout20_50, sout20_51, sout20_52, sout20_53, sout20_54, sout20_55, sout20_56, 
                  sout20_57, sout20_58, sout20_59, sout20_60, sout20_61, sout20_62, sout20_63, sout20_64;
          
    //row21        
    output [21:0] sout21_1, sout21_2, sout21_3, sout21_4, sout21_5, sout21_6, sout21_7, sout21_8,
                  sout21_9, sout21_10, sout21_11, sout21_12, sout21_13, sout21_14, sout21_15, sout21_16,
                  sout21_17, sout21_18, sout21_19, sout21_20, sout21_21, sout21_22, sout21_23, sout21_24, 
                  sout21_25, sout21_26, sout21_27, sout21_28, sout21_29, sout21_30, sout21_31, sout21_32,
                  sout21_33, sout21_34, sout21_35, sout21_36, sout21_37, sout21_38, sout21_39, sout21_40,
                  sout21_41, sout21_42, sout21_43, sout21_44, sout21_45, sout21_46, sout21_47, sout21_48,
                  sout21_49, sout21_50, sout21_51, sout21_52, sout21_53, sout21_54, sout21_55, sout21_56, 
                  sout21_57, sout21_58, sout21_59, sout21_60, sout21_61, sout21_62, sout21_63, sout21_64;
                            
    //row22        
    output [21:0] sout22_1, sout22_2, sout22_3, sout22_4, sout22_5, sout22_6, sout22_7, sout22_8,
                  sout22_9, sout22_10, sout22_11, sout22_12, sout22_13, sout22_14, sout22_15, sout22_16,
                  sout22_17, sout22_18, sout22_19, sout22_20, sout22_21, sout22_22, sout22_23, sout22_24, 
                  sout22_25, sout22_26, sout22_27, sout22_28, sout22_29, sout22_30, sout22_31, sout22_32,
                  sout22_33, sout22_34, sout22_35, sout22_36, sout22_37, sout22_38, sout22_39, sout22_40,
                  sout22_41, sout22_42, sout22_43, sout22_44, sout22_45, sout22_46, sout22_47, sout22_48,
                  sout22_49, sout22_50, sout22_51, sout22_52, sout22_53, sout22_54, sout22_55, sout22_56, 
                  sout22_57, sout22_58, sout22_59, sout22_60, sout22_61, sout22_62, sout22_63, sout22_64;
                         
    //row23       
    output [21:0] sout23_1, sout23_2, sout23_3, sout23_4, sout23_5, sout23_6, sout23_7, sout23_8,
                  sout23_9, sout23_10, sout23_11, sout23_12, sout23_13, sout23_14, sout23_15, sout23_16,
                  sout23_17, sout23_18, sout23_19, sout23_20, sout23_21, sout23_22, sout23_23, sout23_24, 
                  sout23_25, sout23_26, sout23_27, sout23_28, sout23_29, sout23_30, sout23_31, sout23_32,
                  sout23_33, sout23_34, sout23_35, sout23_36, sout23_37, sout23_38, sout23_39, sout23_40,
                  sout23_41, sout23_42, sout23_43, sout23_44, sout23_45, sout23_46, sout23_47, sout23_48,
                  sout23_49, sout23_50, sout23_51, sout23_52, sout23_53, sout23_54, sout23_55, sout23_56, 
                  sout23_57, sout23_58, sout23_59, sout23_60, sout23_61, sout23_62, sout23_63, sout23_64;
                  
    //row24        
    output [21:0] sout24_1, sout24_2, sout24_3, sout24_4, sout24_5, sout24_6, sout24_7, sout24_8,
                  sout24_9, sout24_10, sout24_11, sout24_12, sout24_13, sout24_14, sout24_15, sout24_16,
                  sout24_17, sout24_18, sout24_19, sout24_20, sout24_21, sout24_22, sout24_23, sout24_24, 
                  sout24_25, sout24_26, sout24_27, sout24_28, sout24_29, sout24_30, sout24_31, sout24_32,
                  sout24_33, sout24_34, sout24_35, sout24_36, sout24_37, sout24_38, sout24_39, sout24_40,
                  sout24_41, sout24_42, sout24_43, sout24_44, sout24_45, sout24_46, sout24_47, sout24_48,
                  sout24_49, sout24_50, sout24_51, sout24_52, sout24_53, sout24_54, sout24_55, sout24_56, 
                  sout24_57, sout24_58, sout24_59, sout24_60, sout24_61, sout24_62, sout24_63, sout24_64;
                  
    //row25        
    output [21:0] sout25_1, sout25_2, sout25_3, sout25_4, sout25_5, sout25_6, sout25_7, sout25_8,
                  sout25_9, sout25_10, sout25_11, sout25_12, sout25_13, sout25_14, sout25_15, sout25_16,
                  sout25_17, sout25_18, sout25_19, sout25_20, sout25_21, sout25_22, sout25_23, sout25_24, 
                  sout25_25, sout25_26, sout25_27, sout25_28, sout25_29, sout25_30, sout25_31, sout25_32,
                  sout25_33, sout25_34, sout25_35, sout25_36, sout25_37, sout25_38, sout25_39, sout25_40,
                  sout25_41, sout25_42, sout25_43, sout25_44, sout25_45, sout25_46, sout25_47, sout25_48,
                  sout25_49, sout25_50, sout25_51, sout25_52, sout25_53, sout25_54, sout25_55, sout25_56, 
                  sout25_57, sout25_58, sout25_59, sout25_60, sout25_61, sout25_62, sout25_63, sout25_64;
                 
    //row26        
    output [21:0] sout26_1, sout26_2, sout26_3, sout26_4, sout26_5, sout26_6, sout26_7, sout26_8,
                  sout26_9, sout26_10, sout26_11, sout26_12, sout26_13, sout26_14, sout26_15, sout26_16,
                  sout26_17, sout26_18, sout26_19, sout26_20, sout26_21, sout26_22, sout26_23, sout26_24, 
                  sout26_25, sout26_26, sout26_27, sout26_28, sout26_29, sout26_30, sout26_31, sout26_32,
                  sout26_33, sout26_34, sout26_35, sout26_36, sout26_37, sout26_38, sout26_39, sout26_40,
                  sout26_41, sout26_42, sout26_43, sout26_44, sout26_45, sout26_46, sout26_47, sout26_48,
                  sout26_49, sout26_50, sout26_51, sout26_52, sout26_53, sout26_54, sout26_55, sout26_56, 
                  sout26_57, sout26_58, sout26_59, sout26_60, sout26_61, sout26_62, sout26_63, sout26_64;
                  
    //row27        
    output [21:0] sout27_1, sout27_2, sout27_3, sout27_4, sout27_5, sout27_6, sout27_7, sout27_8,
                  sout27_9, sout27_10, sout27_11, sout27_12, sout27_13, sout27_14, sout27_15, sout27_16,
                  sout27_17, sout27_18, sout27_19, sout27_20, sout27_21, sout27_22, sout27_23, sout27_24, 
                  sout27_25, sout27_26, sout27_27, sout27_28, sout27_29, sout27_30, sout27_31, sout27_32,
                  sout27_33, sout27_34, sout27_35, sout27_36, sout27_37, sout27_38, sout27_39, sout27_40,
                  sout27_41, sout27_42, sout27_43, sout27_44, sout27_45, sout27_46, sout27_47, sout27_48,
                  sout27_49, sout27_50, sout27_51, sout27_52, sout27_53, sout27_54, sout27_55, sout27_56, 
                  sout27_57, sout27_58, sout27_59, sout27_60, sout27_61, sout27_62, sout27_63, sout27_64;
                  
    //row28        
    output [21:0] sout28_1, sout28_2, sout28_3, sout28_4, sout28_5, sout28_6, sout28_7, sout28_8,
                  sout28_9, sout28_10, sout28_11, sout28_12, sout28_13, sout28_14, sout28_15, sout28_16,
                  sout28_17, sout28_18, sout28_19, sout28_20, sout28_21, sout28_22, sout28_23, sout28_24, 
                  sout28_25, sout28_26, sout28_27, sout28_28, sout28_29, sout28_30, sout28_31, sout28_32,
                  sout28_33, sout28_34, sout28_35, sout28_36, sout28_37, sout28_38, sout28_39, sout28_40,
                  sout28_41, sout28_42, sout28_43, sout28_44, sout28_45, sout28_46, sout28_47, sout28_48,
                  sout28_49, sout28_50, sout28_51, sout28_52, sout28_53, sout28_54, sout28_55, sout28_56, 
                  sout28_57, sout28_58, sout28_59, sout28_60, sout28_61, sout28_62, sout28_63, sout28_64;
                  
    //row29       
    output [21:0] sout29_1, sout29_2, sout29_3, sout29_4, sout29_5, sout29_6, sout29_7, sout29_8,
                  sout29_9, sout29_10, sout29_11, sout29_12, sout29_13, sout29_14, sout29_15, sout29_16,
                  sout29_17, sout29_18, sout29_19, sout29_20, sout29_21, sout29_22, sout29_23, sout29_24, 
                  sout29_25, sout29_26, sout29_27, sout29_28, sout29_29, sout29_30, sout29_31, sout29_32,
                  sout29_33, sout29_34, sout29_35, sout29_36, sout29_37, sout29_38, sout29_39, sout29_40,
                  sout29_41, sout29_42, sout29_43, sout29_44, sout29_45, sout29_46, sout29_47, sout29_48,
                  sout29_49, sout29_50, sout29_51, sout29_52, sout29_53, sout29_54, sout29_55, sout29_56, 
                  sout29_57, sout29_58, sout29_59, sout29_60, sout29_61, sout29_62, sout29_63, sout29_64;
                  
    //row30        
    output [21:0] sout30_1, sout30_2, sout30_3, sout30_4, sout30_5, sout30_6, sout30_7, sout30_8,
                  sout30_9, sout30_10, sout30_11, sout30_12, sout30_13, sout30_14, sout30_15, sout30_16,
                  sout30_17, sout30_18, sout30_19, sout30_20, sout30_21, sout30_22, sout30_23, sout30_24, 
                  sout30_25, sout30_26, sout30_27, sout30_28, sout30_29, sout30_30, sout30_31, sout30_32,
                  sout30_33, sout30_34, sout30_35, sout30_36, sout30_37, sout30_38, sout30_39, sout30_40,
                  sout30_41, sout30_42, sout30_43, sout30_44, sout30_45, sout30_46, sout30_47, sout30_48,
                  sout30_49, sout30_50, sout30_51, sout30_52, sout30_53, sout30_54, sout30_55, sout30_56, 
                  sout30_57, sout30_58, sout30_59, sout30_60, sout30_61, sout30_62, sout30_63, sout30_64;
                
    //row31        
    output [21:0] sout31_1, sout31_2, sout31_3, sout31_4, sout31_5, sout31_6, sout31_7, sout31_8,
                  sout31_9, sout31_10, sout31_11, sout31_12, sout31_13, sout31_14, sout31_15, sout31_16,
                  sout31_17, sout31_18, sout31_19, sout31_20, sout31_21, sout31_22, sout31_23, sout31_24, 
                  sout31_25, sout31_26, sout31_27, sout31_28, sout31_29, sout31_30, sout31_31, sout31_32,
                  sout31_33, sout31_34, sout31_35, sout31_36, sout31_37, sout31_38, sout31_39, sout31_40,
                  sout31_41, sout31_42, sout31_43, sout31_44, sout31_45, sout31_46, sout31_47, sout31_48,
                  sout31_49, sout31_50, sout31_51, sout31_52, sout31_53, sout31_54, sout31_55, sout31_56, 
                  sout31_57, sout31_58, sout31_59, sout31_60, sout31_61, sout31_62, sout31_63, sout31_64;
                  
    //row32        
    output [21:0] sout32_1, sout32_2, sout32_3, sout32_4, sout32_5, sout32_6, sout32_7, sout32_8,
                  sout32_9, sout32_10, sout32_11, sout32_12, sout32_13, sout32_14, sout32_15, sout32_16,
                  sout32_17, sout32_18, sout32_19, sout32_20, sout32_21, sout32_22, sout32_23, sout32_24, 
                  sout32_25, sout32_26, sout32_27, sout32_28, sout32_29, sout32_30, sout32_31, sout32_32,
                  sout32_33, sout32_34, sout32_35, sout32_36, sout32_37, sout32_38, sout32_39, sout32_40,
                  sout32_41, sout32_42, sout32_43, sout32_44, sout32_45, sout32_46, sout32_47, sout32_48,
                  sout32_49, sout32_50, sout32_51, sout32_52, sout32_53, sout32_54, sout32_55, sout32_56, 
                  sout32_57, sout32_58, sout32_59, sout32_60, sout32_61, sout32_62, sout32_63, sout32_64;
                  
    //row33        
    output [21:0] sout33_1, sout33_2, sout33_3, sout33_4, sout33_5, sout33_6, sout33_7, sout33_8,
                  sout33_9, sout33_10, sout33_11, sout33_12, sout33_13, sout33_14, sout33_15, sout33_16,
                  sout33_17, sout33_18, sout33_19, sout33_20, sout33_21, sout33_22, sout33_23, sout33_24, 
                  sout33_25, sout33_26, sout33_27, sout33_28, sout33_29, sout33_30, sout33_31, sout33_32,
                  sout33_33, sout33_34, sout33_35, sout33_36, sout33_37, sout33_38, sout33_39, sout33_40,
                  sout33_41, sout33_42, sout33_43, sout33_44, sout33_45, sout33_46, sout33_47, sout33_48,
                  sout33_49, sout33_50, sout33_51, sout33_52, sout33_53, sout33_54, sout33_55, sout33_56, 
                  sout33_57, sout33_58, sout33_59, sout33_60, sout33_61, sout33_62, sout33_63, sout33_64;
                    
                    
    //row34        
    output [21:0] sout34_1, sout34_2, sout34_3, sout34_4, sout34_5, sout34_6, sout34_7, sout34_8,
                  sout34_9, sout34_10, sout34_11, sout34_12, sout34_13, sout34_14, sout34_15, sout34_16,
                  sout34_17, sout34_18, sout34_19, sout34_20, sout34_21, sout34_22, sout34_23, sout34_24, 
                  sout34_25, sout34_26, sout34_27, sout34_28, sout34_29, sout34_30, sout34_31, sout34_32,
                  sout34_33, sout34_34, sout34_35, sout34_36, sout34_37, sout34_38, sout34_39, sout34_40,
                  sout34_41, sout34_42, sout34_43, sout34_44, sout34_45, sout34_46, sout34_47, sout34_48,
                  sout34_49, sout34_50, sout34_51, sout34_52, sout34_53, sout34_54, sout34_55, sout34_56, 
                  sout34_57, sout34_58, sout34_59, sout34_60, sout34_61, sout34_62, sout34_63, sout34_64;
                  
    //row35        
    output [21:0] sout35_1, sout35_2, sout35_3, sout35_4, sout35_5, sout35_6, sout35_7, sout35_8,
                  sout35_9, sout35_10, sout35_11, sout35_12, sout35_13, sout35_14, sout35_15, sout35_16,
                  sout35_17, sout35_18, sout35_19, sout35_20, sout35_21, sout35_22, sout35_23, sout35_24, 
                  sout35_25, sout35_26, sout35_27, sout35_28, sout35_29, sout35_30, sout35_31, sout35_32,
                  sout35_33, sout35_34, sout35_35, sout35_36, sout35_37, sout35_38, sout35_39, sout35_40,
                  sout35_41, sout35_42, sout35_43, sout35_44, sout35_45, sout35_46, sout35_47, sout35_48,
                  sout35_49, sout35_50, sout35_51, sout35_52, sout35_53, sout35_54, sout35_55, sout35_56, 
                  sout35_57, sout35_58, sout35_59, sout35_60, sout35_61, sout35_62, sout35_63, sout35_64;
                  
    //row36        
    output [21:0] sout36_1, sout36_2, sout36_3, sout36_4, sout36_5, sout36_6, sout36_7, sout36_8,
                  sout36_9, sout36_10, sout36_11, sout36_12, sout36_13, sout36_14, sout36_15, sout36_16,
                  sout36_17, sout36_18, sout36_19, sout36_20, sout36_21, sout36_22, sout36_23, sout36_24, 
                  sout36_25, sout36_26, sout36_27, sout36_28, sout36_29, sout36_30, sout36_31, sout36_32,
                  sout36_33, sout36_34, sout36_35, sout36_36, sout36_37, sout36_38, sout36_39, sout36_40,
                  sout36_41, sout36_42, sout36_43, sout36_44, sout36_45, sout36_46, sout36_47, sout36_48,
                  sout36_49, sout36_50, sout36_51, sout36_52, sout36_53, sout36_54, sout36_55, sout36_56, 
                  sout36_57, sout36_58, sout36_59, sout36_60, sout36_61, sout36_62, sout36_63, sout36_64;
                  
    //row37        
    output [21:0] sout37_1, sout37_2, sout37_3, sout37_4, sout37_5, sout37_6, sout37_7, sout37_8,
                  sout37_9, sout37_10, sout37_11, sout37_12, sout37_13, sout37_14, sout37_15, sout37_16,
                  sout37_17, sout37_18, sout37_19, sout37_20, sout37_21, sout37_22, sout37_23, sout37_24, 
                  sout37_25, sout37_26, sout37_27, sout37_28, sout37_29, sout37_30, sout37_31, sout37_32,
                  sout37_33, sout37_34, sout37_35, sout37_36, sout37_37, sout37_38, sout37_39, sout37_40,
                  sout37_41, sout37_42, sout37_43, sout37_44, sout37_45, sout37_46, sout37_47, sout37_48,
                  sout37_49, sout37_50, sout37_51, sout37_52, sout37_53, sout37_54, sout37_55, sout37_56, 
                  sout37_57, sout37_58, sout37_59, sout37_60, sout37_61, sout37_62, sout37_63, sout37_64;
                  
    //row38        
    output [21:0] sout38_1, sout38_2, sout38_3, sout38_4, sout38_5, sout38_6, sout38_7, sout38_8,
                  sout38_9, sout38_10, sout38_11, sout38_12, sout38_13, sout38_14, sout38_15, sout38_16,
                  sout38_17, sout38_18, sout38_19, sout38_20, sout38_21, sout38_22, sout38_23, sout38_24, 
                  sout38_25, sout38_26, sout38_27, sout38_28, sout38_29, sout38_30, sout38_31, sout38_32,
                  sout38_33, sout38_34, sout38_35, sout38_36, sout38_37, sout38_38, sout38_39, sout38_40,
                  sout38_41, sout38_42, sout38_43, sout38_44, sout38_45, sout38_46, sout38_47, sout38_48,
                  sout38_49, sout38_50, sout38_51, sout38_52, sout38_53, sout38_54, sout38_55, sout38_56, 
                  sout38_57, sout38_58, sout38_59, sout38_60, sout38_61, sout38_62, sout38_63, sout38_64;
                  
    //row39        
    output [21:0] sout39_1, sout39_2, sout39_3, sout39_4, sout39_5, sout39_6, sout39_7, sout39_8,
                  sout39_9, sout39_10, sout39_11, sout39_12, sout39_13, sout39_14, sout39_15, sout39_16,
                  sout39_17, sout39_18, sout39_19, sout39_20, sout39_21, sout39_22, sout39_23, sout39_24, 
                  sout39_25, sout39_26, sout39_27, sout39_28, sout39_29, sout39_30, sout39_31, sout39_32,
                  sout39_33, sout39_34, sout39_35, sout39_36, sout39_37, sout39_38, sout39_39, sout39_40,
                  sout39_41, sout39_42, sout39_43, sout39_44, sout39_45, sout39_46, sout39_47, sout39_48,
                  sout39_49, sout39_50, sout39_51, sout39_52, sout39_53, sout39_54, sout39_55, sout39_56, 
                  sout39_57, sout39_58, sout39_59, sout39_60, sout39_61, sout39_62, sout39_63, sout39_64;
                  
    //row40        
    output [21:0] sout40_1, sout40_2, sout40_3, sout40_4, sout40_5, sout40_6, sout40_7, sout40_8,
                  sout40_9, sout40_10, sout40_11, sout40_12, sout40_13, sout40_14, sout40_15, sout40_16,
                  sout40_17, sout40_18, sout40_19, sout40_20, sout40_21, sout40_22, sout40_23, sout40_24, 
                  sout40_25, sout40_26, sout40_27, sout40_28, sout40_29, sout40_30, sout40_31, sout40_32,
                  sout40_33, sout40_34, sout40_35, sout40_36, sout40_37, sout40_38, sout40_39, sout40_40,
                  sout40_41, sout40_42, sout40_43, sout40_44, sout40_45, sout40_46, sout40_47, sout40_48,
                  sout40_49, sout40_50, sout40_51, sout40_52, sout40_53, sout40_54, sout40_55, sout40_56, 
                  sout40_57, sout40_58, sout40_59, sout40_60, sout40_61, sout40_62, sout40_63, sout40_64;
                  
    //row41        
    output [21:0] sout41_1, sout41_2, sout41_3, sout41_4, sout41_5, sout41_6, sout41_7, sout41_8,
                  sout41_9, sout41_10, sout41_11, sout41_12, sout41_13, sout41_14, sout41_15, sout41_16,
                  sout41_17, sout41_18, sout41_19, sout41_20, sout41_21, sout41_22, sout41_23, sout41_24, 
                  sout41_25, sout41_26, sout41_27, sout41_28, sout41_29, sout41_30, sout41_31, sout41_32,
                  sout41_33, sout41_34, sout41_35, sout41_36, sout41_37, sout41_38, sout41_39, sout41_40,
                  sout41_41, sout41_42, sout41_43, sout41_44, sout41_45, sout41_46, sout41_47, sout41_48,
                  sout41_49, sout41_50, sout41_51, sout41_52, sout41_53, sout41_54, sout41_55, sout41_56, 
                  sout41_57, sout41_58, sout41_59, sout41_60, sout41_61, sout41_62, sout41_63, sout41_64;
                  
    //row42        
    output [21:0] sout42_1, sout42_2, sout42_3, sout42_4, sout42_5, sout42_6, sout42_7, sout42_8,
                  sout42_9, sout42_10, sout42_11, sout42_12, sout42_13, sout42_14, sout42_15, sout42_16,
                  sout42_17, sout42_18, sout42_19, sout42_20, sout42_21, sout42_22, sout42_23, sout42_24, 
                  sout42_25, sout42_26, sout42_27, sout42_28, sout42_29, sout42_30, sout42_31, sout42_32,
                  sout42_33, sout42_34, sout42_35, sout42_36, sout42_37, sout42_38, sout42_39, sout42_40,
                  sout42_41, sout42_42, sout42_43, sout42_44, sout42_45, sout42_46, sout42_47, sout42_48,
                  sout42_49, sout42_50, sout42_51, sout42_52, sout42_53, sout42_54, sout42_55, sout42_56, 
                  sout42_57, sout42_58, sout42_59, sout42_60, sout42_61, sout42_62, sout42_63, sout42_64;
                  
    //row43        
    output [21:0] sout43_1, sout43_2, sout43_3, sout43_4, sout43_5, sout43_6, sout43_7, sout43_8,
                  sout43_9, sout43_10, sout43_11, sout43_12, sout43_13, sout43_14, sout43_15, sout43_16,
                  sout43_17, sout43_18, sout43_19, sout43_20, sout43_21, sout43_22, sout43_23, sout43_24, 
                  sout43_25, sout43_26, sout43_27, sout43_28, sout43_29, sout43_30, sout43_31, sout43_32,
                  sout43_33, sout43_34, sout43_35, sout43_36, sout43_37, sout43_38, sout43_39, sout43_40,
                  sout43_41, sout43_42, sout43_43, sout43_44, sout43_45, sout43_46, sout43_47, sout43_48,
                  sout43_49, sout43_50, sout43_51, sout43_52, sout43_53, sout43_54, sout43_55, sout43_56, 
                  sout43_57, sout43_58, sout43_59, sout43_60, sout43_61, sout43_62, sout43_63, sout43_64;
                  
    //row44        
    output [21:0] sout44_1, sout44_2, sout44_3, sout44_4, sout44_5, sout44_6, sout44_7, sout44_8,
                  sout44_9, sout44_10, sout44_11, sout44_12, sout44_13, sout44_14, sout44_15, sout44_16,
                  sout44_17, sout44_18, sout44_19, sout44_20, sout44_21, sout44_22, sout44_23, sout44_24, 
                  sout44_25, sout44_26, sout44_27, sout44_28, sout44_29, sout44_30, sout44_31, sout44_32,
                  sout44_33, sout44_34, sout44_35, sout44_36, sout44_37, sout44_38, sout44_39, sout44_40,
                  sout44_41, sout44_42, sout44_43, sout44_44, sout44_45, sout44_46, sout44_47, sout44_48,
                  sout44_49, sout44_50, sout44_51, sout44_52, sout44_53, sout44_54, sout44_55, sout44_56, 
                  sout44_57, sout44_58, sout44_59, sout44_60, sout44_61, sout44_62, sout44_63, sout44_64;
                  
    //row45        
    output [21:0] sout45_1, sout45_2, sout45_3, sout45_4, sout45_5, sout45_6, sout45_7, sout45_8,
                  sout45_9, sout45_10, sout45_11, sout45_12, sout45_13, sout45_14, sout45_15, sout45_16,
                  sout45_17, sout45_18, sout45_19, sout45_20, sout45_21, sout45_22, sout45_23, sout45_24, 
                  sout45_25, sout45_26, sout45_27, sout45_28, sout45_29, sout45_30, sout45_31, sout45_32,
                  sout45_33, sout45_34, sout45_35, sout45_36, sout45_37, sout45_38, sout45_39, sout45_40,
                  sout45_41, sout45_42, sout45_43, sout45_44, sout45_45, sout45_46, sout45_47, sout45_48,
                  sout45_49, sout45_50, sout45_51, sout45_52, sout45_53, sout45_54, sout45_55, sout45_56, 
                  sout45_57, sout45_58, sout45_59, sout45_60, sout45_61, sout45_62, sout45_63, sout45_64;
                  
    //row46        
    output [21:0] sout46_1, sout46_2, sout46_3, sout46_4, sout46_5, sout46_6, sout46_7, sout46_8,
                  sout46_9, sout46_10, sout46_11, sout46_12, sout46_13, sout46_14, sout46_15, sout46_16,
                  sout46_17, sout46_18, sout46_19, sout46_20, sout46_21, sout46_22, sout46_23, sout46_24, 
                  sout46_25, sout46_26, sout46_27, sout46_28, sout46_29, sout46_30, sout46_31, sout46_32,
                  sout46_33, sout46_34, sout46_35, sout46_36, sout46_37, sout46_38, sout46_39, sout46_40,
                  sout46_41, sout46_42, sout46_43, sout46_44, sout46_45, sout46_46, sout46_47, sout46_48,
                  sout46_49, sout46_50, sout46_51, sout46_52, sout46_53, sout46_54, sout46_55, sout46_56, 
                  sout46_57, sout46_58, sout46_59, sout46_60, sout46_61, sout46_62, sout46_63, sout46_64;
                 
    //row47        
    output [21:0] sout47_1, sout47_2, sout47_3, sout47_4, sout47_5, sout47_6, sout47_7, sout47_8,
                  sout47_9, sout47_10, sout47_11, sout47_12, sout47_13, sout47_14, sout47_15, sout47_16,
                  sout47_17, sout47_18, sout47_19, sout47_20, sout47_21, sout47_22, sout47_23, sout47_24, 
                  sout47_25, sout47_26, sout47_27, sout47_28, sout47_29, sout47_30, sout47_31, sout47_32,
                  sout47_33, sout47_34, sout47_35, sout47_36, sout47_37, sout47_38, sout47_39, sout47_40,
                  sout47_41, sout47_42, sout47_43, sout47_44, sout47_45, sout47_46, sout47_47, sout47_48,
                  sout47_49, sout47_50, sout47_51, sout47_52, sout47_53, sout47_54, sout47_55, sout47_56, 
                  sout47_57, sout47_58, sout47_59, sout47_60, sout47_61, sout47_62, sout47_63, sout47_64;
                  
    //row48        
    output [21:0] sout48_1, sout48_2, sout48_3, sout48_4, sout48_5, sout48_6, sout48_7, sout48_8,
                  sout48_9, sout48_10, sout48_11, sout48_12, sout48_13, sout48_14, sout48_15, sout48_16,
                  sout48_17, sout48_18, sout48_19, sout48_20, sout48_21, sout48_22, sout48_23, sout48_24, 
                  sout48_25, sout48_26, sout48_27, sout48_28, sout48_29, sout48_30, sout48_31, sout48_32,
                  sout48_33, sout48_34, sout48_35, sout48_36, sout48_37, sout48_38, sout48_39, sout48_40,
                  sout48_41, sout48_42, sout48_43, sout48_44, sout48_45, sout48_46, sout48_47, sout48_48,
                  sout48_49, sout48_50, sout48_51, sout48_52, sout48_53, sout48_54, sout48_55, sout48_56, 
                  sout48_57, sout48_58, sout48_59, sout48_60, sout48_61, sout48_62, sout48_63, sout48_64;
                  
    //row49       
    output [21:0] sout49_1, sout49_2, sout49_3, sout49_4, sout49_5, sout49_6, sout49_7, sout49_8,
                  sout49_9, sout49_10, sout49_11, sout49_12, sout49_13, sout49_14, sout49_15, sout49_16,
                  sout49_17, sout49_18, sout49_19, sout49_20, sout49_21, sout49_22, sout49_23, sout49_24, 
                  sout49_25, sout49_26, sout49_27, sout49_28, sout49_29, sout49_30, sout49_31, sout49_32,
                  sout49_33, sout49_34, sout49_35, sout49_36, sout49_37, sout49_38, sout49_39, sout49_40,
                  sout49_41, sout49_42, sout49_43, sout49_44, sout49_45, sout49_46, sout49_47, sout49_48,
                  sout49_49, sout49_50, sout49_51, sout49_52, sout49_53, sout49_54, sout49_55, sout49_56, 
                  sout49_57, sout49_58, sout49_59, sout49_60, sout49_61, sout49_62, sout49_63, sout49_64;
                  
    //row50        
    output [21:0] sout50_1, sout50_2, sout50_3, sout50_4, sout50_5, sout50_6, sout50_7, sout50_8,
                  sout50_9, sout50_10, sout50_11, sout50_12, sout50_13, sout50_14, sout50_15, sout50_16,
                  sout50_17, sout50_18, sout50_19, sout50_20, sout50_21, sout50_22, sout50_23, sout50_24, 
                  sout50_25, sout50_26, sout50_27, sout50_28, sout50_29, sout50_30, sout50_31, sout50_32,
                  sout50_33, sout50_34, sout50_35, sout50_36, sout50_37, sout50_38, sout50_39, sout50_40,
                  sout50_41, sout50_42, sout50_43, sout50_44, sout50_45, sout50_46, sout50_47, sout50_48,
                  sout50_49, sout50_50, sout50_51, sout50_52, sout50_53, sout50_54, sout50_55, sout50_56, 
                  sout50_57, sout50_58, sout50_59, sout50_60, sout50_61, sout50_62, sout50_63, sout50_64;
                  
    //row51        
    output [21:0] sout51_1, sout51_2, sout51_3, sout51_4, sout51_5, sout51_6, sout51_7, sout51_8,
                  sout51_9, sout51_10, sout51_11, sout51_12, sout51_13, sout51_14, sout51_15, sout51_16,
                  sout51_17, sout51_18, sout51_19, sout51_20, sout51_21, sout51_22, sout51_23, sout51_24, 
                  sout51_25, sout51_26, sout51_27, sout51_28, sout51_29, sout51_30, sout51_31, sout51_32,
                  sout51_33, sout51_34, sout51_35, sout51_36, sout51_37, sout51_38, sout51_39, sout51_40,
                  sout51_41, sout51_42, sout51_43, sout51_44, sout51_45, sout51_46, sout51_47, sout51_48,
                  sout51_49, sout51_50, sout51_51, sout51_52, sout51_53, sout51_54, sout51_55, sout51_56, 
                  sout51_57, sout51_58, sout51_59, sout51_60, sout51_61, sout51_62, sout51_63, sout51_64;
                              
    //row52        
    output [21:0] sout52_1, sout52_2, sout52_3, sout52_4, sout52_5, sout52_6, sout52_7, sout52_8,
                  sout52_9, sout52_10, sout52_11, sout52_12, sout52_13, sout52_14, sout52_15, sout52_16,
                  sout52_17, sout52_18, sout52_19, sout52_20, sout52_21, sout52_22, sout52_23, sout52_24, 
                  sout52_25, sout52_26, sout52_27, sout52_28, sout52_29, sout52_30, sout52_31, sout52_32,
                  sout52_33, sout52_34, sout52_35, sout52_36, sout52_37, sout52_38, sout52_39, sout52_40,
                  sout52_41, sout52_42, sout52_43, sout52_44, sout52_45, sout52_46, sout52_47, sout52_48,
                  sout52_49, sout52_50, sout52_51, sout52_52, sout52_53, sout52_54, sout52_55, sout52_56, 
                  sout52_57, sout52_58, sout52_59, sout52_60, sout52_61, sout52_62, sout52_63, sout52_64;
                  
    //row53        
    output [21:0] sout53_1, sout53_2, sout53_3, sout53_4, sout53_5, sout53_6, sout53_7, sout53_8,
                  sout53_9, sout53_10, sout53_11, sout53_12, sout53_13, sout53_14, sout53_15, sout53_16,
                  sout53_17, sout53_18, sout53_19, sout53_20, sout53_21, sout53_22, sout53_23, sout53_24, 
                  sout53_25, sout53_26, sout53_27, sout53_28, sout53_29, sout53_30, sout53_31, sout53_32,
                  sout53_33, sout53_34, sout53_35, sout53_36, sout53_37, sout53_38, sout53_39, sout53_40,
                  sout53_41, sout53_42, sout53_43, sout53_44, sout53_45, sout53_46, sout53_47, sout53_48,
                  sout53_49, sout53_50, sout53_51, sout53_52, sout53_53, sout53_54, sout53_55, sout53_56, 
                  sout53_57, sout53_58, sout53_59, sout53_60, sout53_61, sout53_62, sout53_63, sout53_64;
                  
    //row54        
    output [21:0] sout54_1, sout54_2, sout54_3, sout54_4, sout54_5, sout54_6, sout54_7, sout54_8,
                  sout54_9, sout54_10, sout54_11, sout54_12, sout54_13, sout54_14, sout54_15, sout54_16,
                  sout54_17, sout54_18, sout54_19, sout54_20, sout54_21, sout54_22, sout54_23, sout54_24, 
                  sout54_25, sout54_26, sout54_27, sout54_28, sout54_29, sout54_30, sout54_31, sout54_32,
                  sout54_33, sout54_34, sout54_35, sout54_36, sout54_37, sout54_38, sout54_39, sout54_40,
                  sout54_41, sout54_42, sout54_43, sout54_44, sout54_45, sout54_46, sout54_47, sout54_48,
                  sout54_49, sout54_50, sout54_51, sout54_52, sout54_53, sout54_54, sout54_55, sout54_56, 
                  sout54_57, sout54_58, sout54_59, sout54_60, sout54_61, sout54_62, sout54_63, sout54_64;
                  
    //row55     
    output [21:0] sout55_1, sout55_2, sout55_3, sout55_4, sout55_5, sout55_6, sout55_7, sout55_8,
                  sout55_9, sout55_10, sout55_11, sout55_12, sout55_13, sout55_14, sout55_15, sout55_16,
                  sout55_17, sout55_18, sout55_19, sout55_20, sout55_21, sout55_22, sout55_23, sout55_24, 
                  sout55_25, sout55_26, sout55_27, sout55_28, sout55_29, sout55_30, sout55_31, sout55_32,
                  sout55_33, sout55_34, sout55_35, sout55_36, sout55_37, sout55_38, sout55_39, sout55_40,
                  sout55_41, sout55_42, sout55_43, sout55_44, sout55_45, sout55_46, sout55_47, sout55_48,
                  sout55_49, sout55_50, sout55_51, sout55_52, sout55_53, sout55_54, sout55_55, sout55_56, 
                  sout55_57, sout55_58, sout55_59, sout55_60, sout55_61, sout55_62, sout55_63, sout55_64;
                  
    //row56     
    output [21:0] sout56_1, sout56_2, sout56_3, sout56_4, sout56_5, sout56_6, sout56_7, sout56_8,
                  sout56_9, sout56_10, sout56_11, sout56_12, sout56_13, sout56_14, sout56_15, sout56_16,
                  sout56_17, sout56_18, sout56_19, sout56_20, sout56_21, sout56_22, sout56_23, sout56_24, 
                  sout56_25, sout56_26, sout56_27, sout56_28, sout56_29, sout56_30, sout56_31, sout56_32,
                  sout56_33, sout56_34, sout56_35, sout56_36, sout56_37, sout56_38, sout56_39, sout56_40,
                  sout56_41, sout56_42, sout56_43, sout56_44, sout56_45, sout56_46, sout56_47, sout56_48,
                  sout56_49, sout56_50, sout56_51, sout56_52, sout56_53, sout56_54, sout56_55, sout56_56, 
                  sout56_57, sout56_58, sout56_59, sout56_60, sout56_61, sout56_62, sout56_63, sout56_64;
                  
    //row57     
    output [21:0] sout57_1, sout57_2, sout57_3, sout57_4, sout57_5, sout57_6, sout57_7, sout57_8,
                  sout57_9, sout57_10, sout57_11, sout57_12, sout57_13, sout57_14, sout57_15, sout57_16,
                  sout57_17, sout57_18, sout57_19, sout57_20, sout57_21, sout57_22, sout57_23, sout57_24, 
                  sout57_25, sout57_26, sout57_27, sout57_28, sout57_29, sout57_30, sout57_31, sout57_32,
                  sout57_33, sout57_34, sout57_35, sout57_36, sout57_37, sout57_38, sout57_39, sout57_40,
                  sout57_41, sout57_42, sout57_43, sout57_44, sout57_45, sout57_46, sout57_47, sout57_48,
                  sout57_49, sout57_50, sout57_51, sout57_52, sout57_53, sout57_54, sout57_55, sout57_56, 
                  sout57_57, sout57_58, sout57_59, sout57_60, sout57_61, sout57_62, sout57_63, sout57_64;
                  
    //row58     
    output [21:0] sout58_1, sout58_2, sout58_3, sout58_4, sout58_5, sout58_6, sout58_7, sout58_8,
                  sout58_9, sout58_10, sout58_11, sout58_12, sout58_13, sout58_14, sout58_15, sout58_16,
                  sout58_17, sout58_18, sout58_19, sout58_20, sout58_21, sout58_22, sout58_23, sout58_24, 
                  sout58_25, sout58_26, sout58_27, sout58_28, sout58_29, sout58_30, sout58_31, sout58_32,
                  sout58_33, sout58_34, sout58_35, sout58_36, sout58_37, sout58_38, sout58_39, sout58_40,
                  sout58_41, sout58_42, sout58_43, sout58_44, sout58_45, sout58_46, sout58_47, sout58_48,
                  sout58_49, sout58_50, sout58_51, sout58_52, sout58_53, sout58_54, sout58_55, sout58_56, 
                  sout58_57, sout58_58, sout58_59, sout58_60, sout58_61, sout58_62, sout58_63, sout58_64;
                  
    //row59     
    output [21:0] sout59_1, sout59_2, sout59_3, sout59_4, sout59_5, sout59_6, sout59_7, sout59_8,
                  sout59_9, sout59_10, sout59_11, sout59_12, sout59_13, sout59_14, sout59_15, sout59_16,
                  sout59_17, sout59_18, sout59_19, sout59_20, sout59_21, sout59_22, sout59_23, sout59_24, 
                  sout59_25, sout59_26, sout59_27, sout59_28, sout59_29, sout59_30, sout59_31, sout59_32,
                  sout59_33, sout59_34, sout59_35, sout59_36, sout59_37, sout59_38, sout59_39, sout59_40,
                  sout59_41, sout59_42, sout59_43, sout59_44, sout59_45, sout59_46, sout59_47, sout59_48,
                  sout59_49, sout59_50, sout59_51, sout59_52, sout59_53, sout59_54, sout59_55, sout59_56, 
                  sout59_57, sout59_58, sout59_59, sout59_60, sout59_61, sout59_62, sout59_63, sout59_64;
                  
    //row60     
    output [21:0] sout60_1, sout60_2, sout60_3, sout60_4, sout60_5, sout60_6, sout60_7, sout60_8,
                  sout60_9, sout60_10, sout60_11, sout60_12, sout60_13, sout60_14, sout60_15, sout60_16,
                  sout60_17, sout60_18, sout60_19, sout60_20, sout60_21, sout60_22, sout60_23, sout60_24, 
                  sout60_25, sout60_26, sout60_27, sout60_28, sout60_29, sout60_30, sout60_31, sout60_32,
                  sout60_33, sout60_34, sout60_35, sout60_36, sout60_37, sout60_38, sout60_39, sout60_40,
                  sout60_41, sout60_42, sout60_43, sout60_44, sout60_45, sout60_46, sout60_47, sout60_48,
                  sout60_49, sout60_50, sout60_51, sout60_52, sout60_53, sout60_54, sout60_55, sout60_56, 
                  sout60_57, sout60_58, sout60_59, sout60_60, sout60_61, sout60_62, sout60_63, sout60_64;
                  
    //row61     
    output [21:0] sout61_1, sout61_2, sout61_3, sout61_4, sout61_5, sout61_6, sout61_7, sout61_8,
                  sout61_9, sout61_10, sout61_11, sout61_12, sout61_13, sout61_14, sout61_15, sout61_16,
                  sout61_17, sout61_18, sout61_19, sout61_20, sout61_21, sout61_22, sout61_23, sout61_24, 
                  sout61_25, sout61_26, sout61_27, sout61_28, sout61_29, sout61_30, sout61_31, sout61_32,
                  sout61_33, sout61_34, sout61_35, sout61_36, sout61_37, sout61_38, sout61_39, sout61_40,
                  sout61_41, sout61_42, sout61_43, sout61_44, sout61_45, sout61_46, sout61_47, sout61_48,
                  sout61_49, sout61_50, sout61_51, sout61_52, sout61_53, sout61_54, sout61_55, sout61_56, 
                  sout61_57, sout61_58, sout61_59, sout61_60, sout61_61, sout61_62, sout61_63, sout61_64;
                  
    //row62     
    output [21:0] sout62_1, sout62_2, sout62_3, sout62_4, sout62_5, sout62_6, sout62_7, sout62_8,
                  sout62_9, sout62_10, sout62_11, sout62_12, sout62_13, sout62_14, sout62_15, sout62_16,
                  sout62_17, sout62_18, sout62_19, sout62_20, sout62_21, sout62_22, sout62_23, sout62_24, 
                  sout62_25, sout62_26, sout62_27, sout62_28, sout62_29, sout62_30, sout62_31, sout62_32,
                  sout62_33, sout62_34, sout62_35, sout62_36, sout62_37, sout62_38, sout62_39, sout62_40,
                  sout62_41, sout62_42, sout62_43, sout62_44, sout62_45, sout62_46, sout62_47, sout62_48,
                  sout62_49, sout62_50, sout62_51, sout62_52, sout62_53, sout62_54, sout62_55, sout62_56, 
                  sout62_57, sout62_58, sout62_59, sout62_60, sout62_61, sout62_62, sout62_63, sout62_64;
                  
    //row63     
    output [21:0] sout63_1, sout63_2, sout63_3, sout63_4, sout63_5, sout63_6, sout63_7, sout63_8,
                  sout63_9, sout63_10, sout63_11, sout63_12, sout63_13, sout63_14, sout63_15, sout63_16,
                  sout63_17, sout63_18, sout63_19, sout63_20, sout63_21, sout63_22, sout63_23, sout63_24, 
                  sout63_25, sout63_26, sout63_27, sout63_28, sout63_29, sout63_30, sout63_31, sout63_32,
                  sout63_33, sout63_34, sout63_35, sout63_36, sout63_37, sout63_38, sout63_39, sout63_40,
                  sout63_41, sout63_42, sout63_43, sout63_44, sout63_45, sout63_46, sout63_47, sout63_48,
                  sout63_49, sout63_50, sout63_51, sout63_52, sout63_53, sout63_54, sout63_55, sout63_56, 
                  sout63_57, sout63_58, sout63_59, sout63_60, sout63_61, sout63_62, sout63_63, sout63_64;
                  
    //row64   
    output [21:0] sout64_1, sout64_2, sout64_3, sout64_4, sout64_5, sout64_6, sout64_7, sout64_8,
                  sout64_9, sout64_10, sout64_11, sout64_12, sout64_13, sout64_14, sout64_15, sout64_16,
                  sout64_17, sout64_18, sout64_19, sout64_20, sout64_21, sout64_22, sout64_23, sout64_24, 
                  sout64_25, sout64_26, sout64_27, sout64_28, sout64_29, sout64_30, sout64_31, sout64_32,
                  sout64_33, sout64_34, sout64_35, sout64_36, sout64_37, sout64_38, sout64_39, sout64_40,
                  sout64_41, sout64_42, sout64_43, sout64_44, sout64_45, sout64_46, sout64_47, sout64_48,
                  sout64_49, sout64_50, sout64_51, sout64_52, sout64_53, sout64_54, sout64_55, sout64_56, 
                  sout64_57, sout64_58, sout64_59, sout64_60, sout64_61, sout64_62, sout64_63, sout64_64;
    
      
    //16 4x4 by 16 4x4
    
    //row1
    //mac_array_4x4_11
    wire [7:0] aout14, aout24, aout34, aout44,
               wout41, wout42, wout43, wout44;
                
    //mac_array_4x4_12
    wire [7:0] aout18, aout28, aout38, aout48,
               wout45, wout46, wout47, wout48;
                       
    //mac_array_4x4_13
    wire [7:0] aout1_12, aout2_12, aout3_12, aout4_12,
               wout49, wout4_10, wout4_11, wout4_12;
                
    //mac_array_4x4_14
    wire [7:0] aout1_16, aout2_16, aout3_16, aout4_16,
               wout4_13, wout4_14, wout4_15, wout4_16;
                
    //mac_array_4x4_15
    wire [7:0] aout1_20, aout2_20, aout3_20, aout4_20,
               wout4_17, wout4_18, wout4_19, wout4_20;
                
    //mac_array_4x4_16
    wire [7:0] aout1_24, aout2_24, aout3_24, aout4_24,
               wout4_21, wout4_22, wout4_23, wout4_24;
                
    //mac_array_4x4_17
    wire [7:0] aout1_28, aout2_28, aout3_28, aout4_28,
               wout4_25, wout4_26, wout4_27, wout4_28;
                
    //mac_array_4x4_18
    wire [7:0] aout1_32, aout2_32, aout3_32, aout4_32,
               wout4_29, wout4_30, wout4_31, wout4_32;
                
    //mac_array_4x4_19
    wire [7:0] aout1_36, aout2_36, aout3_36, aout4_36,
               wout4_33, wout4_34, wout4_35, wout4_36;
                            
    //mac_array_4x4_1_10
    wire [7:0] aout1_40, aout2_40, aout3_40, aout4_40,
               wout4_37, wout4_38, wout4_39, wout4_40;
                
    //mac_array_4x4_1_11
    wire [7:0] aout1_44, aout2_44, aout3_44, aout4_44,
               wout4_41, wout4_42, wout4_43, wout4_44;
                
    //mac_array_4x4_1_12
    wire [7:0] aout1_48, aout2_48, aout3_48, aout4_48,
               wout4_45, wout4_46, wout4_47, wout4_48;
                
    //mac_array_4x4_1_13
    wire [7:0] aout1_52, aout2_52, aout3_52, aout4_52,
               wout4_49, wout4_50, wout4_51, wout4_52;
                
    //mac_array_4x4_1_14
    wire [7:0] aout1_56, aout2_56, aout3_56, aout4_56,
               wout4_53, wout4_54, wout4_55, wout4_56;
                
    //mac_array_4x4_1_15
    wire [7:0] aout1_60, aout2_60, aout3_60, aout4_60,
               wout4_57, wout4_58, wout4_59, wout4_60;
                
    //mac_array_4x4_1_16
    wire [7:0] aout1_64, aout2_64, aout3_64, aout4_64,
               wout4_61, wout4_62, wout4_63, wout4_64;
       
   
   
    //row2
    //mac_array_4x4_21
    wire [7:0] aout54, aout64, aout74, aout84,
               wout81, wout82, wout83, wout84;
                
    //mac_array_4x4_22
    wire [7:0] aout58, aout68, aout78, aout88,
               wout85, wout86, wout87, wout88;
                
    //mac_array_4x4_23
    wire [7:0] aout5_12, aout6_12, aout7_12, aout8_12,
               wout89, wout8_10, wout8_11, wout8_12;
                
    //mac_array_4x4_24
    wire [7:0] aout5_16, aout6_16, aout7_16, aout8_16,
               wout8_13, wout8_14, wout8_15, wout8_16;
                
    //mac_array_4x4_25
    wire [7:0] aout5_20, aout6_20, aout7_20, aout8_20,
               wout8_17, wout8_18, wout8_19, wout8_20;
                
    //mac_array_4x4_26
    wire [7:0] aout5_24, aout6_24, aout7_24, aout8_24,
               wout8_21, wout8_22, wout8_23, wout8_24;
                
    //mac_array_4x4_27
    wire [7:0] aout5_28, aout6_28, aout7_28, aout8_28,
               wout8_25, wout8_26, wout8_27, wout8_28;
                
    //mac_array_4x4_28
    wire [7:0] aout5_32, aout6_32, aout7_32, aout8_32,
               wout8_29, wout8_30, wout8_31, wout8_32;
                
    //mac_array_4x4_29
    wire [7:0] aout5_36, aout6_36, aout7_36, aout8_36,
               wout8_33, wout8_34, wout8_35, wout8_36;
                
    //mac_array_4x4_2_10
    wire [7:0] aout5_40, aout6_40, aout7_40, aout8_40,
               wout8_37, wout8_38, wout8_39, wout8_40;
                
    //mac_array_4x4_2_11
    wire [7:0] aout5_44, aout6_44, aout7_44, aout8_44,
               wout8_41, wout8_42, wout8_43, wout8_44;
                
    //mac_array_4x4_2_12
    wire [7:0] aout5_48, aout6_48, aout7_48, aout8_48,
               wout8_45, wout8_46, wout8_47, wout8_48;
                
    //mac_array_4x4_2_13
    wire [7:0] aout5_52, aout6_52, aout7_52, aout8_52,
               wout8_49, wout8_50, wout8_51, wout8_52;
                
    //mac_array_4x4_2_14
    wire [7:0] aout5_56, aout6_56, aout7_56, aout8_56,
               wout8_53, wout8_54, wout8_55, wout8_56;
                
    //mac_array_4x4_2_15
    wire [7:0] aout5_60, aout6_60, aout7_60, aout8_60,
               wout8_57, wout8_58, wout8_59, wout8_60;
                
    //mac_array_4x4_2_16
    wire [7:0] aout5_64, aout6_64, aout7_64, aout8_64,
               wout8_61, wout8_62, wout8_63, wout8_64;
                
                
    
    //row3
    //mac_array_4x4_31
    wire [7:0] aout94, aout10_4, aout11_4, aout12_4,
               wout12_1, wout12_2, wout12_3, wout12_4;
                
    //mac_array_4x4_32
    wire [7:0] aout98, aout10_8, aout11_8, aout12_8,
               wout12_5, wout12_6, wout12_7, wout12_8;
                
    //mac_array_4x4_33
    wire [7:0] aout9_12, aout10_12, aout11_12, aout12_12,
               wout12_9, wout12_10, wout12_11, wout12_12;
                
    //mac_array_4x4_34
    wire [7:0] aout9_16, aout10_16, aout11_16, aout12_16,
               wout12_13, wout12_14, wout12_15, wout12_16;
                
    //mac_array_4x4_35
    wire [7:0] aout9_20, aout10_20, aout11_20, aout12_20,
               wout12_17, wout12_18, wout12_19, wout12_20;
                
    //mac_array_4x4_36
    wire [7:0] aout9_24, aout10_24, aout11_24, aout12_24,
               wout12_21, wout12_22, wout12_23, wout12_24;
                
    //mac_array_4x4_37
    wire [7:0] aout9_28, aout10_28, aout11_28, aout12_28,
               wout12_25, wout12_26, wout12_27, wout12_28;
                
    //mac_array_4x4_38
    wire [7:0] aout9_32, aout10_32, aout11_32, aout12_32,
               wout12_29, wout12_30, wout12_31, wout12_32;
                
    //mac_array_4x4_39
    wire [7:0] aout9_36, aout10_36, aout11_36, aout12_36,
               wout12_33, wout12_34, wout12_35, wout12_36;
                
                
    //mac_array_4x4_3_10
    wire [7:0] aout9_40, aout10_40, aout11_40, aout12_40,
               wout12_37, wout12_38, wout12_39, wout12_40;
                
    //mac_array_4x4_3_11
    wire [7:0] aout9_44, aout10_44, aout11_44, aout12_44,
               wout12_41, wout12_42, wout12_43, wout12_44;
                
    //mac_array_4x4_3_12
    wire [7:0] aout9_48, aout10_48, aout11_48, aout12_48,
               wout12_45, wout12_46, wout12_47, wout12_48;
                
    //mac_array_4x4_3_13
    wire [7:0] aout9_52, aout10_52, aout11_52, aout12_52,
               wout12_49, wout12_50, wout12_51, wout12_52;
                
    //mac_array_4x4_3_14
    wire [7:0] aout9_56, aout10_56, aout11_56, aout12_56,
               wout12_53, wout12_54, wout12_55, wout12_56;
                
    //mac_array_4x4_3_15
    wire [7:0] aout9_60, aout10_60, aout11_60, aout12_60,
               wout12_57, wout12_58, wout12_59, wout12_60;
                
    //mac_array_4x4_3_16
    wire [7:0] aout9_64, aout10_64, aout11_64, aout12_64,
               wout12_61, wout12_62, wout12_63, wout12_64;
       
   
   
    //row4
    //mac_array_4x4_41
    wire [7:0] aout13_4, aout14_4, aout15_4, aout16_4,
               wout16_1, wout16_2, wout16_3, wout16_4;
                
    //mac_array_4x4_42
    wire [7:0] aout13_8, aout14_8, aout15_8, aout16_8,
               wout16_5, wout16_6, wout16_7, wout16_8;
                
    //mac_array_4x4_43
    wire [7:0] aout13_12, aout14_12, aout15_12, aout16_12,
               wout16_9, wout16_10, wout16_11, wout16_12;
                
    //mac_array_4x4_44
    wire [7:0] aout13_16, aout14_16, aout15_16, aout16_16,
               wout16_13, wout16_14, wout16_15, wout16_16;
                
    //mac_array_4x4_45
    wire [7:0] aout13_20, aout14_20, aout15_20, aout16_20,
               wout16_17, wout16_18, wout16_19, wout16_20;
                
    //mac_array_4x4_46
    wire [7:0] aout13_24, aout14_24, aout15_24, aout16_24,
               wout16_21, wout16_22, wout16_23, wout16_24;
                
    //mac_array_4x4_47
    wire [7:0] aout13_28, aout14_28, aout15_28, aout16_28,
               wout16_25, wout16_26, wout16_27, wout16_28;
                
    //mac_array_4x4_48
    wire [7:0] aout13_32, aout14_32, aout15_32, aout16_32,
               wout16_29, wout16_30, wout16_31, wout16_32;
                
    //mac_array_4x4_49
    wire [7:0] aout13_36, aout14_36, aout15_36, aout16_36,
               wout16_33, wout16_34, wout16_35, wout16_36;
                
    //mac_array_4x4_4_10
    wire [7:0] aout13_40, aout14_40, aout15_40, aout16_40,
               wout16_37, wout16_38, wout16_39, wout16_40;
                
    //mac_array_4x4_4_11
    wire [7:0] aout13_44, aout14_44, aout15_44, aout16_44,
               wout16_41, wout16_42, wout16_43, wout16_44;
                
    //mac_array_4x4_4_12
    wire [7:0] aout13_48, aout14_48, aout15_48, aout16_48,
               wout16_45, wout16_46, wout16_47, wout16_48;
                
    //mac_array_4x4_4_13
    wire [7:0] aout13_52, aout14_52, aout15_52, aout16_52,
               wout16_49, wout16_50, wout16_51, wout16_52;
                
    //mac_array_4x4_4_14
    wire [7:0] aout13_56, aout14_56, aout15_56, aout16_56,
               wout16_53, wout16_54, wout16_55, wout16_56;
                
    //mac_array_4x4_4_15
    wire [7:0] aout13_60, aout14_60, aout15_60, aout16_60,
               wout16_57, wout16_58, wout16_59, wout16_60;
                
    //mac_array_4x4_4_16
    wire [7:0] aout13_64, aout14_64, aout15_64, aout16_64,
               wout16_61, wout16_62, wout16_63, wout16_64;
       
       
    //row5
    //mac_array_4x4_51
    wire [7:0] aout17_4, aout18_4, aout19_4, aout20_4,
               wout20_1, wout20_2, wout20_3, wout20_4;
                
    //mac_array_4x4_52
    wire [7:0] aout17_8, aout18_8, aout19_8, aout20_8,
               wout20_5, wout20_6, wout20_7, wout20_8;
                
    //mac_array_4x4_53
    wire [7:0] aout17_12, aout18_12, aout19_12, aout20_12,
               wout20_9, wout20_10, wout20_11, wout20_12;
                
    //mac_array_4x4_54
    wire [7:0] aout17_16, aout18_16, aout19_16, aout20_16,
               wout20_13, wout20_14, wout20_15, wout20_16;
                
    //mac_array_4x4_55
    wire [7:0] aout17_20, aout18_20, aout19_20, aout20_20,
               wout20_17, wout20_18, wout20_19, wout20_20;
                
    //mac_array_4x4_56
    wire [7:0] aout17_24, aout18_24, aout19_24, aout20_24,
               wout20_21, wout20_22, wout20_23, wout20_24;
                
    //mac_array_4x4_57
    wire [7:0] aout17_28, aout18_28, aout19_28, aout20_28,
               wout20_25, wout20_26, wout20_27, wout20_28;
                
    //mac_array_4x4_58
    wire [7:0] aout17_32, aout18_32, aout19_32, aout20_32,
               wout20_29, wout20_30, wout20_31, wout20_32;
                
    //mac_array_4x4_59
    wire [7:0] aout17_36, aout18_36, aout19_36, aout20_36,
               wout20_33, wout20_34, wout20_35, wout20_36;
                
    //mac_array_4x4_5_10
    wire [7:0] aout17_40, aout18_40, aout19_40, aout20_40,
               wout20_37, wout20_38, wout20_39, wout20_40;
                
    //mac_array_4x4_5_11
    wire [7:0] aout17_44, aout18_44, aout19_44, aout20_44,
               wout20_41, wout20_42, wout20_43, wout20_44;
                
    //mac_array_4x4_5_12
    wire [7:0] aout17_48, aout18_48, aout19_48, aout20_48,
               wout20_45, wout20_46, wout20_47, wout20_48;
                
    //mac_array_4x4_5_13
    wire [7:0] aout17_52, aout18_52, aout19_52, aout20_52,
               wout20_49, wout20_50, wout20_51, wout20_52;
                
    //mac_array_4x4_5_14
    wire [7:0] aout17_56, aout18_56, aout19_56, aout20_56,
               wout20_53, wout20_54, wout20_55, wout20_56;
                
    //mac_array_4x4_5_15
    wire [7:0] aout17_60, aout18_60, aout19_60, aout20_60,
               wout20_57, wout20_58, wout20_59, wout20_60;
                
    //mac_array_4x4_5_16
    wire [7:0] aout17_64, aout18_64, aout19_64, aout20_64,
               wout20_61, wout20_62, wout20_63, wout20_64;
               
     
    //row6
    //mac_array_4x4_61
    wire [7:0] aout21_4, aout22_4, aout23_4, aout24_4,
               wout24_1, wout24_2, wout24_3, wout24_4;
                
    //mac_array_4x4_62
    wire [7:0] aout21_8, aout22_8, aout23_8, aout24_8,
               wout24_5, wout24_6, wout24_7, wout24_8;
               
    //mac_array_4x4_63
    wire [7:0] aout21_12, aout22_12, aout23_12, aout24_12,
               wout24_9, wout24_10, wout24_11, wout24_12;
                
    //mac_array_4x4_64
    wire [7:0] aout21_16, aout22_16, aout23_16, aout24_16,
               wout24_13, wout24_14, wout24_15, wout24_16;
                
    //mac_array_4x4_65
    wire [7:0] aout21_20, aout22_20, aout23_20, aout24_20,
               wout24_17, wout24_18, wout24_19, wout24_20;
                
    //mac_array_4x4_66
    wire [7:0] aout21_24, aout22_24, aout23_24, aout24_24,
               wout24_21, wout24_22, wout24_23, wout24_24;
                
    //mac_array_4x4_67
    wire [7:0] aout21_28, aout22_28, aout23_28, aout24_28,
               wout24_25, wout24_26, wout24_27, wout24_28;
                
    //mac_array_4x4_68
    wire [7:0] aout21_32, aout22_32, aout23_32, aout24_32,
               wout24_29, wout24_30, wout24_31, wout24_32;
                
    //mac_array_4x4_69
    wire [7:0] aout21_36, aout22_36, aout23_36, aout24_36,
               wout24_33, wout24_34, wout24_35, wout24_36;
                
    //mac_array_4x4_6_10
    wire [7:0] aout21_40, aout22_40, aout23_40, aout24_40,
               wout24_37, wout24_38, wout24_39, wout24_40;
                
    //mac_array_4x4_6_11
    wire [7:0] aout21_44, aout22_44, aout23_44, aout24_44,
               wout24_41, wout24_42, wout24_43, wout24_44;
                
    //mac_array_4x4_6_12
    wire [7:0] aout21_48, aout22_48, aout23_48, aout24_48,
               wout24_45, wout24_46, wout24_47, wout24_48;
                
    //mac_array_4x4_6_13
    wire [7:0] aout21_52, aout22_52, aout23_52, aout24_52,
               wout24_49, wout24_50, wout24_51, wout24_52;
                
    //mac_array_4x4_6_14
    wire [7:0] aout21_56, aout22_56, aout23_56, aout24_56,
               wout24_53, wout24_54, wout24_55, wout24_56;
                
    //mac_array_4x4_6_15
    wire [7:0] aout21_60, aout22_60, aout23_60, aout24_60,
               wout24_57, wout24_58, wout24_59, wout24_60;
                
    //mac_array_4x4_6_16
    wire [7:0] aout21_64, aout22_64, aout23_64, aout24_64,
               wout24_61, wout24_62, wout24_63, wout24_64;
               
                
    //row7
    //mac_array_4x4_71
    wire [7:0] aout25_4, aout26_4, aout27_4, aout28_4,
               wout28_1, wout28_2, wout28_3, wout28_4;
                
    //mac_array_4x4_72
    wire [7:0] aout25_8, aout26_8, aout27_8, aout28_8,
               wout28_5, wout28_6, wout28_7, wout28_8;
                
    //mac_array_4x4_73
    wire [7:0] aout25_12, aout26_12, aout27_12, aout28_12,
               wout28_9, wout28_10, wout28_11, wout28_12;
                
    //mac_array_4x4_74
    wire [7:0] aout25_16, aout26_16, aout27_16, aout28_16,
               wout28_13, wout28_14, wout28_15, wout28_16;
                
    //mac_array_4x4_75
    wire [7:0] aout25_20, aout26_20, aout27_20, aout28_20,
               wout28_17, wout28_18, wout28_19, wout28_20;
                
    //mac_array_4x4_76
    wire [7:0] aout25_24, aout26_24, aout27_24, aout28_24,
               wout28_21, wout28_22, wout28_23, wout28_24;
                
    //mac_array_4x4_77
    wire [7:0] aout25_28, aout26_28, aout27_28, aout28_28,
               wout28_25, wout28_26, wout28_27, wout28_28;
                
    //mac_array_4x4_78
    wire [7:0] aout25_32, aout26_32, aout27_32, aout28_32,
               wout28_29, wout28_30, wout28_31, wout28_32;
                
    //mac_array_4x4_79
    wire [7:0] aout25_36, aout26_36, aout27_36, aout28_36,
               wout28_33, wout28_34, wout28_35, wout28_36;
                
    //mac_array_4x4_7_10
    wire [7:0] aout25_40, aout26_40, aout27_40, aout28_40,
               wout28_37, wout28_38, wout28_39, wout28_40;
                
    //mac_array_4x4_7_11
    wire [7:0] aout25_44, aout26_44, aout27_44, aout28_44,
               wout28_41, wout28_42, wout28_43, wout28_44;
                
    //mac_array_4x4_7_12
    wire [7:0] aout25_48, aout26_48, aout27_48, aout28_48,
               wout28_45, wout28_46, wout28_47, wout28_48;
                
    //mac_array_4x4_7_13
    wire [7:0] aout25_52, aout26_52, aout27_52, aout28_52,
               wout28_49, wout28_50, wout28_51, wout28_52;
                
    //mac_array_4x4_7_14
    wire [7:0] aout25_56, aout26_56, aout27_56, aout28_56,
               wout28_53, wout28_54, wout28_55, wout28_56;
                
    //mac_array_4x4_7_15
    wire [7:0] aout25_60, aout26_60, aout27_60, aout28_60,
               wout28_57, wout28_58, wout28_59, wout28_60;
                
    //mac_array_4x4_7_16
    wire [7:0] aout25_64, aout26_64, aout27_64, aout28_64,
               wout28_61, wout28_62, wout28_63, wout28_64;
               
              
    //row8
    //mac_array_4x4_81
    wire [7:0] aout29_4, aout30_4, aout31_4, aout32_4,
               wout32_1, wout32_2, wout32_3, wout32_4;
                
    //mac_array_4x4_82
    wire [7:0] aout29_8, aout30_8, aout31_8, aout32_8,
               wout32_5, wout32_6, wout32_7, wout32_8;
                
    //mac_array_4x4_83
    wire [7:0] aout29_12, aout30_12, aout31_12, aout32_12,
               wout32_9, wout32_10, wout32_11, wout32_12;
                
    //mac_array_4x4_84
    wire [7:0] aout29_16, aout30_16, aout31_16, aout32_16,
               wout32_13, wout32_14, wout32_15, wout32_16;
                
    //mac_array_4x4_85
    wire [7:0] aout29_20, aout30_20, aout31_20, aout32_20,
               wout32_17, wout32_18, wout32_19, wout32_20;
                
    //mac_array_4x4_86
    wire [7:0] aout29_24, aout30_24, aout31_24, aout32_24,
               wout32_21, wout32_22, wout32_23, wout32_24;
                
    //mac_array_4x4_87
    wire [7:0] aout29_28, aout30_28, aout31_28, aout32_28,
               wout32_25, wout32_26, wout32_27, wout32_28;
                
    //mac_array_4x4_88
    wire [7:0] aout29_32, aout30_32, aout31_32, aout32_32,
               wout32_29, wout32_30, wout32_31, wout32_32;
                
    //mac_array_4x4_89
    wire [7:0] aout29_36, aout30_36, aout31_36, aout32_36,
               wout32_33, wout32_34, wout32_35, wout32_36;
                
    //mac_array_4x4_8_10
    wire [7:0] aout29_40, aout30_40, aout31_40, aout32_40,
               wout32_37, wout32_38, wout32_39, wout32_40;
                
    //mac_array_4x4_8_11
    wire [7:0] aout29_44, aout30_44, aout31_44, aout32_44,
               wout32_41, wout32_42, wout32_43, wout32_44;
                
    //mac_array_4x4_8_12
    wire [7:0] aout29_48, aout30_48, aout31_48, aout32_48,
               wout32_45, wout32_46, wout32_47, wout32_48;
                
    //mac_array_4x4_8_13
    wire [7:0] aout29_52, aout30_52, aout31_52, aout32_52,
               wout32_49, wout32_50, wout32_51, wout32_52;
                
    //mac_array_4x4_8_14
    wire [7:0] aout29_56, aout30_56, aout31_56, aout32_56,
               wout32_53, wout32_54, wout32_55, wout32_56;
                
    //mac_array_4x4_8_15
    wire [7:0] aout29_60, aout30_60, aout31_60, aout32_60,
               wout32_57, wout32_58, wout32_59, wout32_60;
                
    //mac_array_4x4_8_16
    wire [7:0] aout29_64, aout30_64, aout31_64, aout32_64,
               wout32_61, wout32_62, wout32_63, wout32_64;
       
       
       
    //row9
    //mac_array_4x4_91
    wire [7:0] aout33_4, aout34_4, aout35_4, aout36_4,
               wout36_1, wout36_2, wout36_3, wout36_4;
                
    //mac_array_4x4_92
    wire [7:0] aout33_8, aout34_8, aout35_8, aout36_8,
               wout36_5, wout36_6, wout36_7, wout36_8;
                
    //mac_array_4x4_93
    wire [7:0] aout33_12, aout34_12, aout35_12, aout36_12,
               wout36_9, wout36_10, wout36_11, wout36_12;
                
    //mac_array_4x4_94
    wire [7:0] aout33_16, aout34_16, aout35_16, aout36_16,
               wout36_13, wout36_14, wout36_15, wout36_16;
                
    //mac_array_4x4_95
    wire [7:0] aout33_20, aout34_20, aout35_20, aout36_20,
               wout36_17, wout36_18, wout36_19, wout36_20;
                
    //mac_array_4x4_96
    wire [7:0] aout33_24, aout34_24, aout35_24, aout36_24,
               wout36_21, wout36_22, wout36_23, wout36_24;
                
    //mac_array_4x4_97
    wire [7:0] aout33_28, aout34_28, aout35_28, aout36_28,
               wout36_25, wout36_26, wout36_27, wout36_28;
                
    //mac_array_4x4_98
    wire [7:0] aout33_32, aout34_32, aout35_32, aout36_32,
               wout36_29, wout36_30, wout36_31, wout36_32;
                
    //mac_array_4x4_99
    wire [7:0] aout33_36, aout34_36, aout35_36, aout36_36,
               wout36_33, wout36_34, wout36_35, wout36_36;
                
    //mac_array_4x4_9_10
    wire [7:0] aout33_40, aout34_40, aout35_40, aout36_40,
               wout36_37, wout36_38, wout36_39, wout36_40;
                
    //mac_array_4x4_9_11
    wire [7:0] aout33_44, aout34_44, aout35_44, aout36_44,
               wout36_41, wout36_42, wout36_43, wout36_44;
                
    //mac_array_4x4_9_12
    wire [7:0] aout33_48, aout34_48, aout35_48, aout36_48,
               wout36_45, wout36_46, wout36_47, wout36_48;
                
    //mac_array_4x4_9_13
    wire [7:0] aout33_52, aout34_52, aout35_52, aout36_52,
               wout36_49, wout36_50, wout36_51, wout36_52;
                
    //mac_array_4x4_9_14
    wire [7:0] aout33_56, aout34_56, aout35_56, aout36_56,
               wout36_53, wout36_54, wout36_55, wout36_56;
                
    //mac_array_4x4_9_15
    wire [7:0] aout33_60, aout34_60, aout35_60, aout36_60,
               wout36_57, wout36_58, wout36_59, wout36_60;
                
    //mac_array_4x4_9_16
    wire [7:0] aout33_64, aout34_64, aout35_64, aout36_64,
               wout36_61, wout36_62, wout36_63, wout36_64;
               
  
    //row10
    //mac_array_4x4_10_1
    wire [7:0] aout37_4, aout38_4, aout39_4, aout40_4,
               wout40_1, wout40_2, wout40_3, wout40_4;
                
    //mac_array_4x4_10_2
    wire [7:0] aout37_8, aout38_8, aout39_8, aout40_8,
               wout40_5, wout40_6, wout40_7, wout40_8;
                
    //mac_array_4x4_10_3
    wire [7:0] aout37_12, aout38_12, aout39_12, aout40_12,
               wout40_9, wout40_10, wout40_11, wout40_12;
                
    //mac_array_4x4_10_4
    wire [7:0] aout37_16, aout38_16, aout39_16, aout40_16,
               wout40_13, wout40_14, wout40_15, wout40_16;
                
    //mac_array_4x4_10_5
    wire [7:0] aout37_20, aout38_20, aout39_20, aout40_20,
               wout40_17, wout40_18, wout40_19, wout40_20;
                
    //mac_array_4x4_10_6
    wire [7:0] aout37_24, aout38_24, aout39_24, aout40_24,
               wout40_21, wout40_22, wout40_23, wout40_24;
                
    //mac_array_4x4_10_7
    wire [7:0] aout37_28, aout38_28, aout39_28, aout40_28,
               wout40_25, wout40_26, wout40_27, wout40_28;
                
    //mac_array_4x4_10_8
    wire [7:0] aout37_32, aout38_32, aout39_32, aout40_32,
               wout40_29, wout40_30, wout40_31, wout40_32;
                
    //mac_array_4x4_10_9
    wire [7:0] aout37_36, aout38_36, aout39_36, aout40_36,
               wout40_33, wout40_34, wout40_35, wout40_36;
                
    //mac_array_4x4_10_10
    wire [7:0] aout37_40, aout38_40, aout39_40, aout40_40,
               wout40_37, wout40_38, wout40_39, wout40_40;
                
    //mac_array_4x4_10_11
    wire [7:0] aout37_44, aout38_44, aout39_44, aout40_44,
               wout40_41, wout40_42, wout40_43, wout40_44;
                
    //mac_array_4x4_10_12
    wire [7:0] aout37_48, aout38_48, aout39_48, aout40_48,
               wout40_45, wout40_46, wout40_47, wout40_48;
                
    //mac_array_4x4_10_13
    wire [7:0] aout37_52, aout38_52, aout39_52, aout40_52,
               wout40_49, wout40_50, wout40_51, wout40_52;
                
    //mac_array_4x4_10_14
    wire [7:0] aout37_56, aout38_56, aout39_56, aout40_56,
               wout40_53, wout40_54, wout40_55, wout40_56;
                
    //mac_array_4x4_10_15
    wire [7:0] aout37_60, aout38_60, aout39_60, aout40_60,
               wout40_57, wout40_58, wout40_59, wout40_60;
                
    //mac_array_4x4_10_16
    wire [7:0] aout37_64, aout38_64, aout39_64, aout40_64,
               wout40_61, wout40_62, wout40_63, wout40_64;
               
              
    //row11
    //mac_array_4x4_11_1
    wire [7:0] aout41_4, aout42_4, aout43_4, aout44_4,
               wout44_1, wout44_2, wout44_3, wout44_4;
                
    //mac_array_4x4_11_2
    wire [7:0] aout41_8, aout42_8, aout43_8, aout44_8,
               wout44_5, wout44_6, wout44_7, wout44_8;
                
    //mac_array_4x4_11_3
    wire [7:0] aout41_12, aout42_12, aout43_12, aout44_12,
               wout44_9, wout44_10, wout44_11, wout44_12;
                
    //mac_array_4x4_11_4
    wire [7:0] aout41_16, aout42_16, aout43_16, aout44_16,
               wout44_13, wout44_14, wout44_15, wout44_16;
                
    //mac_array_4x4_11_5
    wire [7:0] aout41_20, aout42_20, aout43_20, aout44_20,
               wout44_17, wout44_18, wout44_19, wout44_20;
                
    //mac_array_4x4_11_6
    wire [7:0] aout41_24, aout42_24, aout43_24, aout44_24,
               wout44_21, wout44_22, wout44_23, wout44_24;
                
    //mac_array_4x4_11_7
    wire [7:0] aout41_28, aout42_28, aout43_28, aout44_28,
               wout44_25, wout44_26, wout44_27, wout44_28;
                
    //mac_array_4x4_11_8
    wire [7:0] aout41_32, aout42_32, aout43_32, aout44_32,
               wout44_29, wout44_30, wout44_31, wout44_32;
                
    //mac_array_4x4_11_9
    wire [7:0] aout41_36, aout42_36, aout43_36, aout44_36,
               wout44_33, wout44_34, wout44_35, wout44_36;
                
    //mac_array_4x4_11_10
    wire [7:0] aout41_40, aout42_40, aout43_40, aout44_40,
               wout44_37, wout44_38, wout44_39, wout44_40;
                
    //mac_array_4x4_11_11
    wire [7:0] aout41_44, aout42_44, aout43_44, aout44_44,
               wout44_41, wout44_42, wout44_43, wout44_44;
                
    //mac_array_4x4_11_12
    wire [7:0] aout41_48, aout42_48, aout43_48, aout44_48,
               wout44_45, wout44_46, wout44_47, wout44_48;
                
    //mac_array_4x4_11_13
    wire [7:0] aout41_52, aout42_52, aout43_52, aout44_52,
               wout44_49, wout44_50, wout44_51, wout44_52;
                
    //mac_array_4x4_11_14
    wire [7:0] aout41_56, aout42_56, aout43_56, aout44_56,
               wout44_53, wout44_54, wout44_55, wout44_56;
                
    //mac_array_4x4_11_15
    wire [7:0] aout41_60, aout42_60, aout43_60, aout44_60,
               wout44_57, wout44_58, wout44_59, wout44_60;
                
    //mac_array_4x4_11_16
    wire [7:0] aout41_64, aout42_64, aout43_64, aout44_64,
               wout44_61, wout44_62, wout44_63, wout44_64;
               
               
    //row12
    //mac_array_4x4_12_1
    wire [7:0] aout45_4, aout46_4, aout47_4, aout48_4,
               wout48_1, wout48_2, wout48_3, wout48_4;
                
    //mac_array_4x4_12_2
    wire [7:0] aout45_8, aout46_8, aout47_8, aout48_8,
               wout48_5, wout48_6, wout48_7, wout48_8;
                
    //mac_array_4x4_12_3
    wire [7:0] aout45_12, aout46_12, aout47_12, aout48_12,
               wout48_9, wout48_10, wout48_11, wout48_12;
                
    //mac_array_4x4_12_4
    wire [7:0] aout45_16, aout46_16, aout47_16, aout48_16,
               wout48_13, wout48_14, wout48_15, wout48_16;
                
    //mac_array_4x4_12_5
    wire [7:0] aout45_20, aout46_20, aout47_20, aout48_20,
               wout48_17, wout48_18, wout48_19, wout48_20;
                
    //mac_array_4x4_12_6
    wire [7:0] aout45_24, aout46_24, aout47_24, aout48_24,
               wout48_21, wout48_22, wout48_23, wout48_24;
                
    //mac_array_4x4_12_7
    wire [7:0] aout45_28, aout46_28, aout47_28, aout48_28,
               wout48_25, wout48_26, wout48_27, wout48_28;
                
    //mac_array_4x4_12_8
    wire [7:0] aout45_32, aout46_32, aout47_32, aout48_32,
               wout48_29, wout48_30, wout48_31, wout48_32;
                
    //mac_array_4x4_12_9
    wire [7:0] aout45_36, aout46_36, aout47_36, aout48_36,
               wout48_33, wout48_34, wout48_35, wout48_36;
                
    //mac_array_4x4_12_10
    wire [7:0] aout45_40, aout46_40, aout47_40, aout48_40,
               wout48_37, wout48_38, wout48_39, wout48_40;
                
    //mac_array_4x4_12_11
    wire [7:0] aout45_44, aout46_44, aout47_44, aout48_44,
               wout48_41, wout48_42, wout48_43, wout48_44;
                
    //mac_array_4x4_12_12
    wire [7:0] aout45_48, aout46_48, aout47_48, aout48_48,
               wout48_45, wout48_46, wout48_47, wout48_48;
                
    //mac_array_4x4_12_13
    wire [7:0] aout45_52, aout46_52, aout47_52, aout48_52,
               wout48_49, wout48_50, wout48_51, wout48_52;
                
    //mac_array_4x4_12_14
    wire [7:0] aout45_56, aout46_56, aout47_56, aout48_56,
               wout48_53, wout48_54, wout48_55, wout48_56;
                
    //mac_array_4x4_12_15
    wire [7:0] aout45_60, aout46_60, aout47_60, aout48_60,
               wout48_57, wout48_58, wout48_59, wout48_60;
                
    //mac_array_4x4_12_16
    wire [7:0] aout45_64, aout46_64, aout47_64, aout48_64,
               wout48_61, wout48_62, wout48_63, wout48_64;
               
               
    //row13
    //mac_array_4x4_13_1
    wire [7:0] aout49_4, aout50_4, aout51_4, aout52_4,
               wout52_1, wout52_2, wout52_3, wout52_4;
                
    //mac_array_4x4_13_2
    wire [7:0] aout49_8, aout50_8, aout51_8, aout52_8,
               wout52_5, wout52_6, wout52_7, wout52_8;
                
    //mac_array_4x4_13_3
    wire [7:0] aout49_12, aout50_12, aout51_12, aout52_12,
               wout52_9, wout52_10, wout52_11, wout52_12;
                
    //mac_array_4x4_13_4
    wire [7:0] aout49_16, aout50_16, aout51_16, aout52_16,
               wout52_13, wout52_14, wout52_15, wout52_16;
                
    //mac_array_4x4_13_5
    wire [7:0] aout49_20, aout50_20, aout51_20, aout52_20,
               wout52_17, wout52_18, wout52_19, wout52_20;
                
    //mac_array_4x4_13_6
    wire [7:0] aout49_24, aout50_24, aout51_24, aout52_24,
               wout52_21, wout52_22, wout52_23, wout52_24;
                
    //mac_array_4x4_13_7
    wire [7:0] aout49_28, aout50_28, aout51_28, aout52_28,
               wout52_25, wout52_26, wout52_27, wout52_28;
                
    //mac_array_4x4_13_8
    wire [7:0] aout49_32, aout50_32, aout51_32, aout52_32,
               wout52_29, wout52_30, wout52_31, wout52_32;
                
    //mac_array_4x4_13_9
    wire [7:0] aout49_36, aout50_36, aout51_36, aout52_36,
               wout52_33, wout52_34, wout52_35, wout52_36;
                
    //mac_array_4x4_13_10
    wire [7:0] aout49_40, aout50_40, aout51_40, aout52_40,
               wout52_37, wout52_38, wout52_39, wout52_40;
                
    //mac_array_4x4_13_11
    wire [7:0] aout49_44, aout50_44, aout51_44, aout52_44,
               wout52_41, wout52_42, wout52_43, wout52_44;
                
    //mac_array_4x4_13_12
    wire [7:0] aout49_48, aout50_48, aout51_48, aout52_48,
               wout52_45, wout52_46, wout52_47, wout52_48;
                
    //mac_array_4x4_13_13
    wire [7:0] aout49_52, aout50_52, aout51_52, aout52_52,
               wout52_49, wout52_50, wout52_51, wout52_52;
                
    //mac_array_4x4_13_14
    wire [7:0] aout49_56, aout50_56, aout51_56, aout52_56,
               wout52_53, wout52_54, wout52_55, wout52_56;
                
    //mac_array_4x4_13_15
    wire [7:0] aout49_60, aout50_60, aout51_60, aout52_60,
               wout52_57, wout52_58, wout52_59, wout52_60;
                
    //mac_array_4x4_13_16
    wire [7:0] aout49_64, aout50_64, aout51_64, aout52_64,
               wout52_61, wout52_62, wout52_63, wout52_64;
               
               
    //row14
    //mac_array_4x4_14_1
    wire [7:0] aout53_4, aout54_4, aout55_4, aout56_4,
               wout56_1, wout56_2, wout56_3, wout56_4;
                
    //mac_array_4x4_14_2
    wire [7:0] aout53_8, aout54_8, aout55_8, aout56_8,
               wout56_5, wout56_6, wout56_7, wout56_8;
                
    //mac_array_4x4_14_3
    wire [7:0] aout53_12, aout54_12, aout55_12, aout56_12,
               wout56_9, wout56_10, wout56_11, wout56_12;
                
    //mac_array_4x4_14_4
    wire [7:0] aout53_16, aout54_16, aout55_16, aout56_16,
               wout56_13, wout56_14, wout56_15, wout56_16;
                
    //mac_array_4x4_14_5
    wire [7:0] aout53_20, aout54_20, aout55_20, aout56_20,
               wout56_17, wout56_18, wout56_19, wout56_20;
                
    //mac_array_4x4_14_6
    wire [7:0] aout53_24, aout54_24, aout55_24, aout56_24,
               wout56_21, wout56_22, wout56_23, wout56_24;
                
    //mac_array_4x4_14_7
    wire [7:0] aout53_28, aout54_28, aout55_28, aout56_28,
               wout56_25, wout56_26, wout56_27, wout56_28;
                
    //mac_array_4x4_14_8
    wire [7:0] aout53_32, aout54_32, aout55_32, aout56_32,
               wout56_29, wout56_30, wout56_31, wout56_32;
                
    //mac_array_4x4_14_9
    wire [7:0] aout53_36, aout54_36, aout55_36, aout56_36,
               wout56_33, wout56_34, wout56_35, wout56_36;
                
    //mac_array_4x4_14_10
    wire [7:0] aout53_40, aout54_40, aout55_40, aout56_40,
               wout56_37, wout56_38, wout56_39, wout56_40;
                
    //mac_array_4x4_14_11
    wire [7:0] aout53_44, aout54_44, aout55_44, aout56_44,
               wout56_41, wout56_42, wout56_43, wout56_44;
                
    //mac_array_4x4_14_12
    wire [7:0] aout53_48, aout54_48, aout55_48, aout56_48,
               wout56_45, wout56_46, wout56_47, wout56_48;
                
    //mac_array_4x4_14_13
    wire [7:0] aout53_52, aout54_52, aout55_52, aout56_52,
               wout56_49, wout56_50, wout56_51, wout56_52;
                
    //mac_array_4x4_14_14
    wire [7:0] aout53_56, aout54_56, aout55_56, aout56_56,
               wout56_53, wout56_54, wout56_55, wout56_56;
                
    //mac_array_4x4_14_15
    wire [7:0] aout53_60, aout54_60, aout55_60, aout56_60,
               wout56_57, wout56_58, wout56_59, wout56_60;
                
    //mac_array_4x4_14_16
    wire [7:0] aout53_64, aout54_64, aout55_64, aout56_64,
               wout56_61, wout56_62, wout56_63, wout56_64;
               
               
    //row15
    //mac_array_4x4_15_1
    wire [7:0] aout57_4, aout58_4, aout59_4, aout60_4,
               wout60_1, wout60_2, wout60_3, wout60_4;
                
    //mac_array_4x4_15_2
    wire [7:0] aout57_8, aout58_8, aout59_8, aout60_8,
               wout60_5, wout60_6, wout60_7, wout60_8;
                
    //mac_array_4x4_15_3
    wire [7:0] aout57_12, aout58_12, aout59_12, aout60_12,
               wout60_9, wout60_10, wout60_11, wout60_12;
                
    //mac_array_4x4_15_4
    wire [7:0] aout57_16, aout58_16, aout59_16, aout60_16,
               wout60_13, wout60_14, wout60_15, wout60_16;
                
    //mac_array_4x4_15_5
    wire [7:0] aout57_20, aout58_20, aout59_20, aout60_20,
               wout60_17, wout60_18, wout60_19, wout60_20;
                
    //mac_array_4x4_15_6
    wire [7:0] aout57_24, aout58_24, aout59_24, aout60_24,
               wout60_21, wout60_22, wout60_23, wout60_24;
                
    //mac_array_4x4_15_7
    wire [7:0] aout57_28, aout58_28, aout59_28, aout60_28,
               wout60_25, wout60_26, wout60_27, wout60_28;
                
    //mac_array_4x4_15_8
    wire [7:0] aout57_32, aout58_32, aout59_32, aout60_32,
               wout60_29, wout60_30, wout60_31, wout60_32;
                
    //mac_array_4x4_15_9
    wire [7:0] aout57_36, aout58_36, aout59_36, aout60_36,
               wout60_33, wout60_34, wout60_35, wout60_36;
                
    //mac_array_4x4_15_10
    wire [7:0] aout57_40, aout58_40, aout59_40, aout60_40,
               wout60_37, wout60_38, wout60_39, wout60_40;
                
    //mac_array_4x4_15_11
    wire [7:0] aout57_44, aout58_44, aout59_44, aout60_44,
               wout60_41, wout60_42, wout60_43, wout60_44;
                
    //mac_array_4x4_15_12
    wire [7:0] aout57_48, aout58_48, aout59_48, aout60_48,
               wout60_45, wout60_46, wout60_47, wout60_48;
                
    //mac_array_4x4_15_13
    wire [7:0] aout57_52, aout58_52, aout59_52, aout60_52,
               wout60_49, wout60_50, wout60_51, wout60_52;
                
    //mac_array_4x4_15_14
    wire [7:0] aout57_56, aout58_56, aout59_56, aout60_56,
               wout60_53, wout60_54, wout60_55, wout60_56;
                
    //mac_array_4x4_15_15
    wire [7:0] aout57_60, aout58_60, aout59_60, aout60_60,
               wout60_57, wout60_58, wout60_59, wout60_60;
                
    //mac_array_4x4_15_16
    wire [7:0] aout57_64, aout58_64, aout59_64, aout60_64,
               wout60_61, wout60_62, wout60_63, wout60_64;
       
    
    //row16
    //mac_array_4x4_16_1
    wire [7:0] aout61_4, aout62_4, aout63_4, aout64_4,
               wout64_1, wout64_2, wout64_3, wout64_4;
                
    //mac_array_4x4_16_2
    wire [7:0] aout61_8, aout62_8, aout63_8, aout64_8,
               wout64_5, wout64_6, wout64_7, wout64_8;
                
    //mac_array_4x4_16_3
    wire [7:0] aout61_12, aout62_12, aout63_12, aout64_12,
               wout64_9, wout64_10, wout64_11, wout64_12;
                
    //mac_array_4x4_16_4
    wire [7:0] aout61_16, aout62_16, aout63_16, aout64_16,
               wout64_13, wout64_14, wout64_15, wout64_16;
                
    //mac_array_4x4_16_5
    wire [7:0] aout61_20, aout62_20, aout63_20, aout64_20,
               wout64_17, wout64_18, wout64_19, wout64_20;
                
    //mac_array_4x4_16_6
    wire [7:0] aout61_24, aout62_24, aout63_24, aout64_24,
               wout64_21, wout64_22, wout64_23, wout64_24;
                
    //mac_array_4x4_16_7
    wire [7:0] aout61_28, aout62_28, aout63_28, aout64_28,
               wout64_25, wout64_26, wout64_27, wout64_28;
                
    //mac_array_4x4_16_8
    wire [7:0] aout61_32, aout62_32, aout63_32, aout64_32,
               wout64_29, wout64_30, wout64_31, wout64_32;
                
    //mac_array_4x4_16_9
    wire [7:0] aout61_36, aout62_36, aout63_36, aout64_36,
               wout64_33, wout64_34, wout64_35, wout64_36;
                
    //mac_array_4x4_16_10
    wire [7:0] aout61_40, aout62_40, aout63_40, aout64_40,
               wout64_37, wout64_38, wout64_39, wout64_40;
                
    //mac_array_4x4_16_11
    wire [7:0] aout61_44, aout62_44, aout63_44, aout64_44,
               wout64_41, wout64_42, wout64_43, wout64_44;
                
    //mac_array_4x4_16_12
    wire [7:0] aout61_48, aout62_48, aout63_48, aout64_48,
               wout64_45, wout64_46, wout64_47, wout64_48;
                
    //mac_array_4x4_16_13
    wire [7:0] aout61_52, aout62_52, aout63_52, aout64_52,
               wout64_49, wout64_50, wout64_51, wout64_52;
                
    //mac_array_4x4_16_14
    wire [7:0] aout61_56, aout62_56, aout63_56, aout64_56,
               wout64_53, wout64_54, wout64_55, wout64_56;
                
    //mac_array_4x4_16_15
    wire [7:0] aout61_60, aout62_60, aout63_60, aout64_60,
               wout64_57, wout64_58, wout64_59, wout64_60;
                
    //mac_array_4x4_16_16
    wire [7:0] aout61_64, aout62_64, aout63_64, aout64_64,
               wout64_61, wout64_62, wout64_63, wout64_64;
       
       
       
    //row1
    mac_array_4x4 mac_array_4x4_11 (.clk(clk), .rst(rst),
                    .ain1(ain1), .ain2(ain2), .ain3(ain3), .ain4(ain4),
                    .win1(win1), .win2(win2), .win3(win3), .win4(win4),
                    .aout1(aout14), .aout2(aout24), .aout3(aout34), .aout4(aout44),
                    .wout1(wout41), .wout2(wout42), .wout3(wout43), .wout4(wout44),
                    .sout11(sout11), .sout12(sout12), .sout13(sout13), .sout14(sout14),
                    .sout21(sout21), .sout22(sout22), .sout23(sout23), .sout24(sout24),
                    .sout31(sout31), .sout32(sout32), .sout33(sout33), .sout34(sout34),
                    .sout41(sout41), .sout42(sout42), .sout43(sout43), .sout44(sout44)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_12 (.clk(clk), .rst(rst),
                    .ain1(aout14), .ain2(aout24), .ain3(aout34), .ain4(aout44),
                    .win1(win5), .win2(win6), .win3(win7), .win4(win8),
                    .aout1(aout18), .aout2(aout28), .aout3(aout38), .aout4(aout48),
                    .wout1(wout45), .wout2(wout46), .wout3(wout47), .wout4(wout48),
                    .sout11(sout15), .sout12(sout16), .sout13(sout17), .sout14(sout18),
                    .sout21(sout25), .sout22(sout26), .sout23(sout27), .sout24(sout28),
                    .sout31(sout35), .sout32(sout36), .sout33(sout37), .sout34(sout38),
                    .sout41(sout45), .sout42(sout46), .sout43(sout47), .sout44(sout48)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_13 (.clk(clk), .rst(rst),
                    .ain1(aout18), .ain2(aout28), .ain3(aout38), .ain4(aout48),
                    .win1(win9), .win2(win10), .win3(win11), .win4(win12),
                    .aout1(aout1_12), .aout2(aout2_12), .aout3(aout3_12), .aout4(aout4_12),
                    .wout1(wout49), .wout2(wout4_10), .wout3(wout4_11), .wout4(wout4_12),
                    .sout11(sout19), .sout12(sout1_10), .sout13(sout1_11), .sout14(sout1_12),
                    .sout21(sout29), .sout22(sout2_10), .sout23(sout2_11), .sout24(sout2_12),
                    .sout31(sout39), .sout32(sout3_10), .sout33(sout3_11), .sout34(sout3_12),
                    .sout41(sout49), .sout42(sout4_10), .sout43(sout4_11), .sout44(sout4_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14 (.clk(clk), .rst(rst),
                    .ain1(aout1_12), .ain2(aout2_12), .ain3(aout3_12), .ain4(aout4_12),
                    .win1(win13), .win2(win14), .win3(win15), .win4(win16),
                    .aout1(aout1_16), .aout2(aout2_16), .aout3(aout3_16), .aout4(aout4_16),
                    .wout1(wout4_13), .wout2(wout4_14), .wout3(wout4_15), .wout4(wout4_16),
                    .sout11(sout1_13), .sout12(sout1_14), .sout13(sout1_15), .sout14(sout1_16),
                    .sout21(sout2_13), .sout22(sout2_14), .sout23(sout2_15), .sout24(sout2_16),
                    .sout31(sout3_13), .sout32(sout3_14), .sout33(sout3_15), .sout34(sout3_16),
                    .sout41(sout4_13), .sout42(sout4_14), .sout43(sout4_15), .sout44(sout4_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15 (.clk(clk), .rst(rst),
                    .ain1(aout1_16), .ain2(aout2_16), .ain3(aout3_16), .ain4(aout4_16),
                    .win1(win17), .win2(win18), .win3(win19), .win4(win20),
                    .aout1(aout1_20), .aout2(aout2_20), .aout3(aout3_20), .aout4(aout4_20),
                    .wout1(wout4_17), .wout2(wout4_18), .wout3(wout4_19), .wout4(wout4_20),
                    .sout11(sout1_17), .sout12(sout1_18), .sout13(sout1_19), .sout14(sout1_20),
                    .sout21(sout2_17), .sout22(sout2_18), .sout23(sout2_19), .sout24(sout2_20),
                    .sout31(sout3_17), .sout32(sout3_18), .sout33(sout3_19), .sout34(sout3_20),
                    .sout41(sout4_17), .sout42(sout4_18), .sout43(sout4_19), .sout44(sout4_20)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16 (.clk(clk), .rst(rst),
                    .ain1(aout1_20), .ain2(aout2_20), .ain3(aout3_20), .ain4(aout4_20),
                    .win1(win21), .win2(win22), .win3(win23), .win4(win24),
                    .aout1(aout1_24), .aout2(aout2_24), .aout3(aout3_24), .aout4(aout4_24),
                    .wout1(wout4_21), .wout2(wout4_22), .wout3(wout4_23), .wout4(wout4_24),
                    .sout11(sout1_21), .sout12(sout1_22), .sout13(sout1_23), .sout14(sout1_24),
                    .sout21(sout2_21), .sout22(sout2_22), .sout23(sout2_23), .sout24(sout2_24),
                    .sout31(sout3_21), .sout32(sout3_22), .sout33(sout3_23), .sout34(sout3_24),
                    .sout41(sout4_21), .sout42(sout4_22), .sout43(sout4_23), .sout44(sout4_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_17 (.clk(clk), .rst(rst),
                    .ain1(aout1_24), .ain2(aout2_24), .ain3(aout3_24), .ain4(aout4_24),
                    .win1(win25), .win2(win26), .win3(win27), .win4(win28),
                    .aout1(aout1_28), .aout2(aout2_28), .aout3(aout3_28), .aout4(aout4_28),
                    .wout1(wout4_25), .wout2(wout4_26), .wout3(wout4_27), .wout4(wout4_28),
                    .sout11(sout1_25), .sout12(sout1_26), .sout13(sout1_27), .sout14(sout1_28),
                    .sout21(sout2_25), .sout22(sout2_26), .sout23(sout2_27), .sout24(sout2_28),
                    .sout31(sout3_25), .sout32(sout3_26), .sout33(sout3_27), .sout34(sout3_28),
                    .sout41(sout4_25), .sout42(sout4_26), .sout43(sout4_27), .sout44(sout4_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_18 (.clk(clk), .rst(rst),
                    .ain1(aout1_28), .ain2(aout2_28), .ain3(aout3_28), .ain4(aout4_28),
                    .win1(win29), .win2(win30), .win3(win31), .win4(win32),
                    .aout1(aout1_32), .aout2(aout2_32), .aout3(aout3_32), .aout4(aout4_32),
                    .wout1(wout4_29), .wout2(wout4_30), .wout3(wout4_31), .wout4(wout4_32),
                    .sout11(sout1_29), .sout12(sout1_30), .sout13(sout1_31), .sout14(sout1_32),
                    .sout21(sout2_29), .sout22(sout2_30), .sout23(sout2_31), .sout24(sout2_32),
                    .sout31(sout3_29), .sout32(sout3_30), .sout33(sout3_31), .sout34(sout3_32),
                    .sout41(sout4_29), .sout42(sout4_30), .sout43(sout4_31), .sout44(sout4_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_19 (.clk(clk), .rst(rst),
                    .ain1(aout1_32), .ain2(aout2_32), .ain3(aout3_32), .ain4(aout4_32),
                    .win1(win33), .win2(win34), .win3(win35), .win4(win36),
                    .aout1(aout1_36), .aout2(aout2_36), .aout3(aout3_36), .aout4(aout4_36),
                    .wout1(wout4_33), .wout2(wout4_34), .wout3(wout4_35), .wout4(wout4_36),
                    .sout11(sout1_33), .sout12(sout1_34), .sout13(sout1_35), .sout14(sout1_36),
                    .sout21(sout2_33), .sout22(sout2_34), .sout23(sout2_35), .sout24(sout2_36),
                    .sout31(sout3_33), .sout32(sout3_34), .sout33(sout3_35), .sout34(sout3_36),
                    .sout41(sout4_33), .sout42(sout4_34), .sout43(sout4_35), .sout44(sout4_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_1_10 (.clk(clk), .rst(rst),
                    .ain1(aout1_36), .ain2(aout2_36), .ain3(aout3_36), .ain4(aout4_36),
                    .win1(win37), .win2(win38), .win3(win39), .win4(win40),
                    .aout1(aout1_40), .aout2(aout2_40), .aout3(aout3_40), .aout4(aout4_40),
                    .wout1(wout4_37), .wout2(wout4_38), .wout3(wout4_39), .wout4(wout4_40),
                    .sout11(sout1_37), .sout12(sout1_38), .sout13(sout1_39), .sout14(sout1_40),
                    .sout21(sout2_37), .sout22(sout2_38), .sout23(sout2_39), .sout24(sout2_40),
                    .sout31(sout3_37), .sout32(sout3_38), .sout33(sout3_39), .sout34(sout3_40),
                    .sout41(sout4_37), .sout42(sout4_38), .sout43(sout4_39), .sout44(sout4_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_1_11 (.clk(clk), .rst(rst),
                    .ain1(aout1_40), .ain2(aout2_40), .ain3(aout3_40), .ain4(aout4_40),
                    .win1(win41), .win2(win42), .win3(win43), .win4(win44),
                    .aout1(aout1_44), .aout2(aout2_44), .aout3(aout3_44), .aout4(aout4_44),
                    .wout1(wout4_41), .wout2(wout4_42), .wout3(wout4_43), .wout4(wout4_44),
                    .sout11(sout1_41), .sout12(sout1_42), .sout13(sout1_43), .sout14(sout1_44),
                    .sout21(sout2_41), .sout22(sout2_42), .sout23(sout2_43), .sout24(sout2_44),
                    .sout31(sout3_41), .sout32(sout3_42), .sout33(sout3_43), .sout34(sout3_44),
                    .sout41(sout4_41), .sout42(sout4_42), .sout43(sout4_43), .sout44(sout4_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_1_12 (.clk(clk), .rst(rst),
                    .ain1(aout1_44), .ain2(aout2_44), .ain3(aout3_44), .ain4(aout4_44),
                    .win1(win45), .win2(win46), .win3(win47), .win4(win48),
                    .aout1(aout1_48), .aout2(aout2_48), .aout3(aout3_48), .aout4(aout4_48),
                    .wout1(wout4_45), .wout2(wout4_46), .wout3(wout4_47), .wout4(wout4_48),
                    .sout11(sout1_45), .sout12(sout1_46), .sout13(sout1_47), .sout14(sout1_48),
                    .sout21(sout2_45), .sout22(sout2_46), .sout23(sout2_47), .sout24(sout2_48),
                    .sout31(sout3_45), .sout32(sout3_46), .sout33(sout3_47), .sout34(sout3_48),
                    .sout41(sout4_45), .sout42(sout4_46), .sout43(sout4_47), .sout44(sout4_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_1_13 (.clk(clk), .rst(rst),
                    .ain1(aout1_48), .ain2(aout2_48), .ain3(aout3_48), .ain4(aout4_48),
                    .win1(win49), .win2(win50), .win3(win51), .win4(win52),
                    .aout1(aout1_52), .aout2(aout2_52), .aout3(aout3_52), .aout4(aout4_52),
                    .wout1(wout4_49), .wout2(wout4_50), .wout3(wout4_51), .wout4(wout4_52),
                    .sout11(sout1_49), .sout12(sout1_50), .sout13(sout1_51), .sout14(sout1_52),
                    .sout21(sout2_49), .sout22(sout2_50), .sout23(sout2_51), .sout24(sout2_52),
                    .sout31(sout3_49), .sout32(sout3_50), .sout33(sout3_51), .sout34(sout3_52),
                    .sout41(sout4_49), .sout42(sout4_50), .sout43(sout4_51), .sout44(sout4_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_1_14 (.clk(clk), .rst(rst),
                    .ain1(aout1_52), .ain2(aout2_52), .ain3(aout3_52), .ain4(aout4_52),
                    .win1(win53), .win2(win54), .win3(win55), .win4(win56),
                    .aout1(aout1_56), .aout2(aout2_56), .aout3(aout3_56), .aout4(aout4_56),
                    .wout1(wout4_53), .wout2(wout4_54), .wout3(wout4_55), .wout4(wout4_56),
                    .sout11(sout1_53), .sout12(sout1_54), .sout13(sout1_55), .sout14(sout1_56),
                    .sout21(sout2_53), .sout22(sout2_54), .sout23(sout2_55), .sout24(sout2_56),
                    .sout31(sout3_53), .sout32(sout3_54), .sout33(sout3_55), .sout34(sout3_56),
                    .sout41(sout4_53), .sout42(sout4_54), .sout43(sout4_55), .sout44(sout4_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_1_15 (.clk(clk), .rst(rst),
                    .ain1(aout1_56), .ain2(aout2_56), .ain3(aout3_56), .ain4(aout4_56),
                    .win1(win57), .win2(win58), .win3(win59), .win4(win60),
                    .aout1(aout1_60), .aout2(aout2_60), .aout3(aout3_60), .aout4(aout4_60),
                    .wout1(wout4_57), .wout2(wout4_58), .wout3(wout4_59), .wout4(wout4_60),
                    .sout11(sout1_57), .sout12(sout1_58), .sout13(sout1_59), .sout14(sout1_60),
                    .sout21(sout2_57), .sout22(sout2_58), .sout23(sout2_59), .sout24(sout2_60),
                    .sout31(sout3_57), .sout32(sout3_58), .sout33(sout3_59), .sout34(sout3_60),
                    .sout41(sout4_57), .sout42(sout4_58), .sout43(sout4_59), .sout44(sout4_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_1_16 (.clk(clk), .rst(rst),
                    .ain1(aout1_60), .ain2(aout2_60), .ain3(aout3_60), .ain4(aout4_60),
                    .win1(win61), .win2(win62), .win3(win63), .win4(win64),
                    .aout1(aout1_64), .aout2(aout2_64), .aout3(aout3_64), .aout4(aout4_64),
                    .wout1(wout4_61), .wout2(wout4_62), .wout3(wout4_63), .wout4(wout4_64),
                    .sout11(sout1_61), .sout12(sout1_62), .sout13(sout1_63), .sout14(sout1_64),
                    .sout21(sout2_61), .sout22(sout2_62), .sout23(sout2_63), .sout24(sout2_64),
                    .sout31(sout3_61), .sout32(sout3_62), .sout33(sout3_63), .sout34(sout3_64),
                    .sout41(sout4_61), .sout42(sout4_62), .sout43(sout4_63), .sout44(sout4_64)
                    ); //4x4 MAC array
    
    
    
    //row2 
    mac_array_4x4 mac_array_4x4_21 (.clk(clk), .rst(rst),
                    .ain1(ain5), .ain2(ain6), .ain3(ain7), .ain4(ain8),
                    .win1(wout41), .win2(wout42), .win3(wout43), .win4(wout44),
                    .aout1(aout54), .aout2(aout64), .aout3(aout74), .aout4(aout84),
                    .wout1(wout81), .wout2(wout82), .wout3(wout83), .wout4(wout84),
                    .sout11(sout51), .sout12(sout52), .sout13(sout53), .sout14(sout54),
                    .sout21(sout61), .sout22(sout62), .sout23(sout63), .sout24(sout64),
                    .sout31(sout71), .sout32(sout72), .sout33(sout73), .sout34(sout74),
                    .sout41(sout81), .sout42(sout82), .sout43(sout83), .sout44(sout84)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_22 (.clk(clk), .rst(rst),
                    .ain1(aout54), .ain2(aout64), .ain3(aout74), .ain4(aout84),
                    .win1(wout45), .win2(wout46), .win3(wout47), .win4(wout48),
                    .aout1(aout58), .aout2(aout68), .aout3(aout78), .aout4(aout88),
                    .wout1(wout85), .wout2(wout86), .wout3(wout87), .wout4(wout88),
                    .sout11(sout55), .sout12(sout56), .sout13(sout57), .sout14(sout58),
                    .sout21(sout65), .sout22(sout66), .sout23(sout67), .sout24(sout68),
                    .sout31(sout75), .sout32(sout76), .sout33(sout77), .sout34(sout78),
                    .sout41(sout85), .sout42(sout86), .sout43(sout87), .sout44(sout88)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_23 (.clk(clk), .rst(rst),
                    .ain1(aout58), .ain2(aout68), .ain3(aout78), .ain4(aout88),
                    .win1(wout49), .win2(wout4_10), .win3(wout4_11), .win4(wout4_12),
                    .aout1(aout5_12), .aout2(aout6_12), .aout3(aout7_12), .aout4(aout8_12),
                    .wout1(wout89), .wout2(wout8_10), .wout3(wout8_11), .wout4(wout8_12),
                    .sout11(sout59), .sout12(sout5_10), .sout13(sout5_11), .sout14(sout5_12),
                    .sout21(sout69), .sout22(sout6_10), .sout23(sout6_11), .sout24(sout6_12),
                    .sout31(sout79), .sout32(sout7_10), .sout33(sout7_11), .sout34(sout7_12),
                    .sout41(sout89), .sout42(sout8_10), .sout43(sout8_11), .sout44(sout8_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_24 (.clk(clk), .rst(rst),
                    .ain1(aout5_12), .ain2(aout6_12), .ain3(aout7_12), .ain4(aout8_12),
                    .win1(wout4_13), .win2(wout4_14), .win3(wout4_15), .win4(wout4_16),
                    .aout1(aout5_16), .aout2(aout6_16), .aout3(aout7_16), .aout4(aout8_16),
                    .wout1(wout8_13), .wout2(wout8_14), .wout3(wout8_15), .wout4(wout8_16),
                    .sout11(sout5_13), .sout12(sout5_14), .sout13(sout5_15), .sout14(sout5_16),
                    .sout21(sout6_13), .sout22(sout6_14), .sout23(sout6_15), .sout24(sout6_16),
                    .sout31(sout7_13), .sout32(sout7_14), .sout33(sout7_15), .sout34(sout7_16),
                    .sout41(sout8_13), .sout42(sout8_14), .sout43(sout8_15), .sout44(sout8_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_25 (.clk(clk), .rst(rst),
                    .ain1(aout5_16), .ain2(aout6_16), .ain3(aout7_16), .ain4(aout8_16),
                    .win1(wout4_17), .win2(wout4_18), .win3(wout4_19), .win4(wout4_20),
                    .aout1(aout5_20), .aout2(aout6_20), .aout3(aout7_20), .aout4(aout8_20),
                    .wout1(wout8_17), .wout2(wout8_18), .wout3(wout8_19), .wout4(wout8_20),
                    .sout11(sout5_17), .sout12(sout5_18), .sout13(sout5_19), .sout14(sout5_20),
                    .sout21(sout6_17), .sout22(sout6_18), .sout23(sout6_19), .sout24(sout6_20),
                    .sout31(sout7_17), .sout32(sout7_18), .sout33(sout7_19), .sout34(sout7_20),
                    .sout41(sout8_17), .sout42(sout8_18), .sout43(sout8_19), .sout44(sout8_20)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_26 (.clk(clk), .rst(rst),
                    .ain1(aout5_20), .ain2(aout6_20), .ain3(aout7_20), .ain4(aout8_20),
                    .win1(wout4_21), .win2(wout4_22), .win3(wout4_23), .win4(wout4_24),
                    .aout1(aout5_24), .aout2(aout6_24), .aout3(aout7_24), .aout4(aout8_24),
                    .wout1(wout8_21), .wout2(wout8_22), .wout3(wout8_23), .wout4(wout8_24),
                    .sout11(sout5_21), .sout12(sout5_22), .sout13(sout5_23), .sout14(sout5_24),
                    .sout21(sout6_21), .sout22(sout6_22), .sout23(sout6_23), .sout24(sout6_24),
                    .sout31(sout7_21), .sout32(sout7_22), .sout33(sout7_23), .sout34(sout7_24),
                    .sout41(sout8_21), .sout42(sout8_22), .sout43(sout8_23), .sout44(sout8_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_27 (.clk(clk), .rst(rst),
                    .ain1(aout5_24), .ain2(aout6_24), .ain3(aout7_24), .ain4(aout8_24),
                    .win1(wout4_25), .win2(wout4_26), .win3(wout4_27), .win4(wout4_28),
                    .aout1(aout5_28), .aout2(aout6_28), .aout3(aout7_28), .aout4(aout8_28),
                    .wout1(wout8_25), .wout2(wout8_26), .wout3(wout8_27), .wout4(wout8_28),
                    .sout11(sout5_25), .sout12(sout5_26), .sout13(sout5_27), .sout14(sout5_28),
                    .sout21(sout6_25), .sout22(sout6_26), .sout23(sout6_27), .sout24(sout6_28),
                    .sout31(sout7_25), .sout32(sout7_26), .sout33(sout7_27), .sout34(sout7_28),
                    .sout41(sout8_25), .sout42(sout8_26), .sout43(sout8_27), .sout44(sout8_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_28 (.clk(clk), .rst(rst),
                    .ain1(aout5_28), .ain2(aout6_28), .ain3(aout7_28), .ain4(aout8_28),
                    .win1(wout4_29), .win2(wout4_30), .win3(wout4_31), .win4(wout4_32),
                    .aout1(aout5_32), .aout2(aout6_32), .aout3(aout7_32), .aout4(aout8_32),
                    .wout1(wout8_29), .wout2(wout8_30), .wout3(wout8_31), .wout4(wout8_32),
                    .sout11(sout5_29), .sout12(sout5_30), .sout13(sout5_31), .sout14(sout5_32),
                    .sout21(sout6_29), .sout22(sout6_30), .sout23(sout6_31), .sout24(sout6_32),
                    .sout31(sout7_29), .sout32(sout7_30), .sout33(sout7_31), .sout34(sout7_32),
                    .sout41(sout8_29), .sout42(sout8_30), .sout43(sout8_31), .sout44(sout8_32)
                    ); //4x4 MAC array
                                  
    mac_array_4x4 mac_array_4x4_29 (.clk(clk), .rst(rst),
                    .ain1(aout5_32), .ain2(aout6_32), .ain3(aout7_32), .ain4(aout8_32),
                    .win1(wout4_33), .win2(wout4_34), .win3(wout4_35), .win4(wout4_36),
                    .aout1(aout5_36), .aout2(aout6_36), .aout3(aout7_36), .aout4(aout8_36),
                    .wout1(wout8_33), .wout2(wout8_34), .wout3(wout8_35), .wout4(wout8_36),
                    .sout11(sout5_33), .sout12(sout5_34), .sout13(sout5_35), .sout14(sout5_36),
                    .sout21(sout6_33), .sout22(sout6_34), .sout23(sout6_35), .sout24(sout6_36),
                    .sout31(sout7_33), .sout32(sout7_34), .sout33(sout7_35), .sout34(sout7_36),
                    .sout41(sout8_33), .sout42(sout8_34), .sout43(sout8_35), .sout44(sout8_36)
                    ); //4x4 MAC array
        
                
    mac_array_4x4 mac_array_4x4_2_10 (.clk(clk), .rst(rst),
                    .ain1(aout5_36), .ain2(aout6_36), .ain3(aout7_36), .ain4(aout8_36),
                    .win1(wout4_37), .win2(wout4_38), .win3(wout4_39), .win4(wout4_40),
                    .aout1(aout5_40), .aout2(aout6_40), .aout3(aout7_40), .aout4(aout8_40),
                    .wout1(wout8_37), .wout2(wout8_38), .wout3(wout8_39), .wout4(wout8_40),
                    .sout11(sout5_37), .sout12(sout5_38), .sout13(sout5_39), .sout14(sout5_40),
                    .sout21(sout6_37), .sout22(sout6_38), .sout23(sout6_39), .sout24(sout6_40),
                    .sout31(sout7_37), .sout32(sout7_38), .sout33(sout7_39), .sout34(sout7_40),
                    .sout41(sout8_37), .sout42(sout8_38), .sout43(sout8_39), .sout44(sout8_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_2_11 (.clk(clk), .rst(rst),
                    .ain1(aout5_40), .ain2(aout6_40), .ain3(aout7_40), .ain4(aout8_40),
                    .win1(wout4_41), .win2(wout4_42), .win3(wout4_43), .win4(wout4_44),
                    .aout1(aout5_44), .aout2(aout6_44), .aout3(aout7_44), .aout4(aout8_44),
                    .wout1(wout8_41), .wout2(wout8_42), .wout3(wout8_43), .wout4(wout8_44),
                    .sout11(sout5_41), .sout12(sout5_42), .sout13(sout5_43), .sout14(sout5_44),
                    .sout21(sout6_41), .sout22(sout6_42), .sout23(sout6_43), .sout24(sout6_44),
                    .sout31(sout7_41), .sout32(sout7_42), .sout33(sout7_43), .sout34(sout7_44),
                    .sout41(sout8_41), .sout42(sout8_42), .sout43(sout8_43), .sout44(sout8_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_2_12 (.clk(clk), .rst(rst),
                    .ain1(aout5_44), .ain2(aout6_44), .ain3(aout7_44), .ain4(aout8_44),
                    .win1(wout4_45), .win2(wout4_46), .win3(wout4_47), .win4(wout4_48),
                    .aout1(aout5_48), .aout2(aout6_48), .aout3(aout7_48), .aout4(aout8_48),
                    .wout1(wout8_45), .wout2(wout8_46), .wout3(wout8_47), .wout4(wout8_48),
                    .sout11(sout5_45), .sout12(sout5_46), .sout13(sout5_47), .sout14(sout5_48),
                    .sout21(sout6_45), .sout22(sout6_46), .sout23(sout6_47), .sout24(sout6_48),
                    .sout31(sout7_45), .sout32(sout7_46), .sout33(sout7_47), .sout34(sout7_48),
                    .sout41(sout8_45), .sout42(sout8_46), .sout43(sout8_47), .sout44(sout8_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_2_13 (.clk(clk), .rst(rst),
                    .ain1(aout5_48), .ain2(aout6_48), .ain3(aout7_48), .ain4(aout8_48),
                    .win1(wout4_49), .win2(wout4_50), .win3(wout4_51), .win4(wout4_52),
                    .aout1(aout5_52), .aout2(aout6_52), .aout3(aout7_52), .aout4(aout8_52),
                    .wout1(wout8_49), .wout2(wout8_50), .wout3(wout8_51), .wout4(wout8_52),
                    .sout11(sout5_49), .sout12(sout5_50), .sout13(sout5_51), .sout14(sout5_52),
                    .sout21(sout6_49), .sout22(sout6_50), .sout23(sout6_51), .sout24(sout6_52),
                    .sout31(sout7_49), .sout32(sout7_50), .sout33(sout7_51), .sout34(sout7_52),
                    .sout41(sout8_49), .sout42(sout8_50), .sout43(sout8_51), .sout44(sout8_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_2_14 (.clk(clk), .rst(rst),
                    .ain1(aout5_52), .ain2(aout6_52), .ain3(aout7_52), .ain4(aout8_52),
                    .win1(wout4_53), .win2(wout4_54), .win3(wout4_55), .win4(wout4_56),
                    .aout1(aout5_56), .aout2(aout6_56), .aout3(aout7_56), .aout4(aout8_56),
                    .wout1(wout8_53), .wout2(wout8_54), .wout3(wout8_55), .wout4(wout8_56),
                    .sout11(sout5_53), .sout12(sout5_54), .sout13(sout5_55), .sout14(sout5_56),
                    .sout21(sout6_53), .sout22(sout6_54), .sout23(sout6_55), .sout24(sout6_56),
                    .sout31(sout7_53), .sout32(sout7_54), .sout33(sout7_55), .sout34(sout7_56),
                    .sout41(sout8_53), .sout42(sout8_54), .sout43(sout8_55), .sout44(sout8_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_2_15 (.clk(clk), .rst(rst),
                    .ain1(aout5_56), .ain2(aout6_56), .ain3(aout7_56), .ain4(aout8_56),
                    .win1(wout4_57), .win2(wout4_58), .win3(wout4_59), .win4(wout4_60),
                    .aout1(aout5_60), .aout2(aout6_60), .aout3(aout7_60), .aout4(aout8_60),
                    .wout1(wout8_57), .wout2(wout8_58), .wout3(wout8_59), .wout4(wout8_60),
                    .sout11(sout5_57), .sout12(sout5_58), .sout13(sout5_59), .sout14(sout5_60),
                    .sout21(sout6_57), .sout22(sout6_58), .sout23(sout6_59), .sout24(sout6_60),
                    .sout31(sout7_57), .sout32(sout7_58), .sout33(sout7_59), .sout34(sout7_60),
                    .sout41(sout8_57), .sout42(sout8_58), .sout43(sout8_59), .sout44(sout8_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_2_16 (.clk(clk), .rst(rst),
                    .ain1(aout5_60), .ain2(aout6_60), .ain3(aout7_60), .ain4(aout8_60),
                    .win1(wout4_61), .win2(wout4_62), .win3(wout4_63), .win4(wout4_64),
                    .aout1(aout5_64), .aout2(aout6_64), .aout3(aout7_64), .aout4(aout8_64),
                    .wout1(wout8_61), .wout2(wout8_62), .wout3(wout8_63), .wout4(wout8_64),
                    .sout11(sout5_61), .sout12(sout5_62), .sout13(sout5_63), .sout14(sout5_64),
                    .sout21(sout6_61), .sout22(sout6_62), .sout23(sout6_63), .sout24(sout6_64),
                    .sout31(sout7_61), .sout32(sout7_62), .sout33(sout7_63), .sout34(sout7_64),
                    .sout41(sout8_61), .sout42(sout8_62), .sout43(sout8_63), .sout44(sout8_64)
                    ); //4x4 MAC array
          
           
                    
    //row 3
    mac_array_4x4 mac_array_4x4_31 (.clk(clk), .rst(rst),
                    .ain1(ain9), .ain2(ain10), .ain3(ain11), .ain4(ain12),
                    .win1(wout81), .win2(wout82), .win3(wout83), .win4(wout84),
                    .aout1(aout94), .aout2(aout10_4), .aout3(aout11_4), .aout4(aout12_4),
                    .wout1(wout12_1), .wout2(wout12_2), .wout3(wout12_3), .wout4(wout12_4),
                    .sout11(sout91), .sout12(sout92), .sout13(sout93), .sout14(sout94),
                    .sout21(sout10_1), .sout22(sout10_2), .sout23(sout10_3), .sout24(sout10_4),
                    .sout31(sout11_1), .sout32(sout11_2), .sout33(sout11_3), .sout34(sout11_4),
                    .sout41(sout12_1), .sout42(sout12_2), .sout43(sout12_3), .sout44(sout12_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_32 (.clk(clk), .rst(rst),
                    .ain1(aout94), .ain2(aout10_4), .ain3(aout11_4), .ain4(aout12_4),
                    .win1(wout85), .win2(wout86), .win3(wout87), .win4(wout88),
                    .aout1(aout98), .aout2(aout10_8), .aout3(aout11_8), .aout4(aout12_8),
                    .wout1(wout12_5), .wout2(wout12_6), .wout3(wout12_7), .wout4(wout12_8),
                    .sout11(sout95), .sout12(sout96), .sout13(sout97), .sout14(sout98),
                    .sout21(sout10_5), .sout22(sout10_6), .sout23(sout10_7), .sout24(sout10_8),
                    .sout31(sout11_5), .sout32(sout11_6), .sout33(sout11_7), .sout34(sout11_8),
                    .sout41(sout12_5), .sout42(sout12_6), .sout43(sout12_7), .sout44(sout12_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_33 (.clk(clk), .rst(rst),
                    .ain1(aout98), .ain2(aout10_8), .ain3(aout11_8), .ain4(aout12_8),
                    .win1(wout89), .win2(wout8_10), .win3(wout8_11), .win4(wout8_12),
                    .aout1(aout9_12), .aout2(aout10_12), .aout3(aout11_12), .aout4(aout12_12),
                    .wout1(wout12_9), .wout2(wout12_10), .wout3(wout12_11), .wout4(wout12_12),
                    .sout11(sout99), .sout12(sout9_10), .sout13(sout9_11), .sout14(sout9_12),
                    .sout21(sout10_9), .sout22(sout10_10), .sout23(sout10_11), .sout24(sout10_12),
                    .sout31(sout11_9), .sout32(sout11_10), .sout33(sout11_11), .sout34(sout11_12),
                    .sout41(sout12_9), .sout42(sout12_10), .sout43(sout12_11), .sout44(sout12_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_34 (.clk(clk), .rst(rst),
                    .ain1(aout9_12), .ain2(aout10_12), .ain3(aout11_12), .ain4(aout12_12),
                    .win1(wout8_13), .win2(wout8_14), .win3(wout8_15), .win4(wout8_16),
                    .aout1(aout9_16), .aout2(aout10_16), .aout3(aout11_16), .aout4(aout12_16),
                    .wout1(wout12_13), .wout2(wout12_14), .wout3(wout12_15), .wout4(wout12_16),
                    .sout11(sout9_13), .sout12(sout9_14), .sout13(sout9_15), .sout14(sout9_16),
                    .sout21(sout10_13), .sout22(sout10_14), .sout23(sout10_15), .sout24(sout10_16),
                    .sout31(sout11_13), .sout32(sout11_14), .sout33(sout11_15), .sout34(sout11_16),
                    .sout41(sout12_13), .sout42(sout12_14), .sout43(sout12_15), .sout44(sout12_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_35 (.clk(clk), .rst(rst),
                    .ain1(aout9_16), .ain2(aout10_16), .ain3(aout11_16), .ain4(aout12_16),
                    .win1(wout8_17), .win2(wout8_18), .win3(wout8_19), .win4(wout8_20),
                    .aout1(aout9_20), .aout2(aout10_20), .aout3(aout11_20), .aout4(aout12_20),
                    .wout1(wout12_17), .wout2(wout12_18), .wout3(wout12_19), .wout4(wout12_20),
                    .sout11(sout9_17), .sout12(sout9_18), .sout13(sout9_19), .sout14(sout9_20),
                    .sout21(sout10_17), .sout22(sout10_18), .sout23(sout10_19), .sout24(sout10_20),
                    .sout31(sout11_17), .sout32(sout11_18), .sout33(sout11_19), .sout34(sout11_20),
                    .sout41(sout12_17), .sout42(sout12_18), .sout43(sout12_19), .sout44(sout12_20)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_36 (.clk(clk), .rst(rst),
                    .ain1(aout9_20), .ain2(aout10_20), .ain3(aout11_20), .ain4(aout12_20),
                    .win1(wout8_21), .win2(wout8_22), .win3(wout8_23), .win4(wout8_24),
                    .aout1(aout9_24), .aout2(aout10_24), .aout3(aout11_24), .aout4(aout12_24),
                    .wout1(wout12_21), .wout2(wout12_22), .wout3(wout12_23), .wout4(wout12_24),
                    .sout11(sout9_21), .sout12(sout9_22), .sout13(sout9_23), .sout14(sout9_24),
                    .sout21(sout10_21), .sout22(sout10_22), .sout23(sout10_23), .sout24(sout10_24),
                    .sout31(sout11_21), .sout32(sout11_22), .sout33(sout11_23), .sout34(sout11_24),
                    .sout41(sout12_21), .sout42(sout12_22), .sout43(sout12_23), .sout44(sout12_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_37 (.clk(clk), .rst(rst),
                    .ain1(aout9_24), .ain2(aout10_24), .ain3(aout11_24), .ain4(aout12_24),
                    .win1(wout8_25), .win2(wout8_26), .win3(wout8_27), .win4(wout8_28),
                    .aout1(aout9_28), .aout2(aout10_28), .aout3(aout11_28), .aout4(aout12_28),
                    .wout1(wout12_25), .wout2(wout12_26), .wout3(wout12_27), .wout4(wout12_28),
                    .sout11(sout9_25), .sout12(sout9_26), .sout13(sout9_27), .sout14(sout9_28),
                    .sout21(sout10_25), .sout22(sout10_26), .sout23(sout10_27), .sout24(sout10_28),
                    .sout31(sout11_25), .sout32(sout11_26), .sout33(sout11_27), .sout34(sout11_28),
                    .sout41(sout12_25), .sout42(sout12_26), .sout43(sout12_27), .sout44(sout12_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_38 (.clk(clk), .rst(rst),
                    .ain1(aout9_28), .ain2(aout10_28), .ain3(aout11_28), .ain4(aout12_28),
                    .win1(wout8_29), .win2(wout8_30), .win3(wout8_31), .win4(wout8_32),
                    .aout1(aout9_32), .aout2(aout10_32), .aout3(aout11_32), .aout4(aout12_32),
                    .wout1(wout12_29), .wout2(wout12_30), .wout3(wout12_31), .wout4(wout12_32),
                    .sout11(sout9_29), .sout12(sout9_30), .sout13(sout9_31), .sout14(sout9_32),
                    .sout21(sout10_29), .sout22(sout10_30), .sout23(sout10_31), .sout24(sout10_32),
                    .sout31(sout11_29), .sout32(sout11_30), .sout33(sout11_31), .sout34(sout11_32),
                    .sout41(sout12_29), .sout42(sout12_30), .sout43(sout12_31), .sout44(sout12_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_39 (.clk(clk), .rst(rst),
                    .ain1(aout9_32), .ain2(aout10_32), .ain3(aout11_32), .ain4(aout12_32),
                    .win1(wout8_33), .win2(wout8_34), .win3(wout8_35), .win4(wout8_36),
                    .aout1(aout9_36), .aout2(aout10_36), .aout3(aout11_36), .aout4(aout12_36),
                    .wout1(wout12_33), .wout2(wout12_34), .wout3(wout12_35), .wout4(wout12_36),
                    .sout11(sout9_33), .sout12(sout9_34), .sout13(sout9_35), .sout14(sout9_36),
                    .sout21(sout10_33), .sout22(sout10_34), .sout23(sout10_35), .sout24(sout10_36),
                    .sout31(sout11_33), .sout32(sout11_34), .sout33(sout11_35), .sout34(sout11_36),
                    .sout41(sout12_33), .sout42(sout12_34), .sout43(sout12_35), .sout44(sout12_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_3_10 (.clk(clk), .rst(rst),
                    .ain1(aout9_36), .ain2(aout10_36), .ain3(aout11_36), .ain4(aout12_36),
                    .win1(wout8_37), .win2(wout8_38), .win3(wout8_39), .win4(wout8_40),
                    .aout1(aout9_40), .aout2(aout10_40), .aout3(aout11_40), .aout4(aout12_40),
                    .wout1(wout12_37), .wout2(wout12_38), .wout3(wout12_39), .wout4(wout12_40),
                    .sout11(sout9_37), .sout12(sout9_38), .sout13(sout9_39), .sout14(sout9_40),
                    .sout21(sout10_37), .sout22(sout10_38), .sout23(sout10_39), .sout24(sout10_40),
                    .sout31(sout11_37), .sout32(sout11_38), .sout33(sout11_39), .sout34(sout11_40),
                    .sout41(sout12_37), .sout42(sout12_38), .sout43(sout12_39), .sout44(sout12_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_3_11 (.clk(clk), .rst(rst),
                    .ain1(aout9_40), .ain2(aout10_40), .ain3(aout11_40), .ain4(aout12_40),
                    .win1(wout8_41), .win2(wout8_42), .win3(wout8_43), .win4(wout8_44),
                    .aout1(aout9_44), .aout2(aout10_44), .aout3(aout11_44), .aout4(aout12_44),
                    .wout1(wout12_41), .wout2(wout12_42), .wout3(wout12_43), .wout4(wout12_44),
                    .sout11(sout9_41), .sout12(sout9_42), .sout13(sout9_43), .sout14(sout9_44),
                    .sout21(sout10_41), .sout22(sout10_42), .sout23(sout10_43), .sout24(sout10_44),
                    .sout31(sout11_41), .sout32(sout11_42), .sout33(sout11_43), .sout34(sout11_44),
                    .sout41(sout12_41), .sout42(sout12_42), .sout43(sout12_43), .sout44(sout12_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_3_12 (.clk(clk), .rst(rst),
                    .ain1(aout9_44), .ain2(aout10_44), .ain3(aout11_44), .ain4(aout12_44),
                    .win1(wout8_45), .win2(wout8_46), .win3(wout8_47), .win4(wout8_48),
                    .aout1(aout9_48), .aout2(aout10_48), .aout3(aout11_48), .aout4(aout12_48),
                    .wout1(wout12_45), .wout2(wout12_46), .wout3(wout12_47), .wout4(wout12_48),
                    .sout11(sout9_45), .sout12(sout9_46), .sout13(sout9_47), .sout14(sout9_48),
                    .sout21(sout10_45), .sout22(sout10_46), .sout23(sout10_47), .sout24(sout10_48),
                    .sout31(sout11_45), .sout32(sout11_46), .sout33(sout11_47), .sout34(sout11_48),
                    .sout41(sout12_45), .sout42(sout12_46), .sout43(sout12_47), .sout44(sout12_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_3_13 (.clk(clk), .rst(rst),
                    .ain1(aout9_48), .ain2(aout10_48), .ain3(aout11_48), .ain4(aout12_48),
                    .win1(wout8_49), .win2(wout8_50), .win3(wout8_51), .win4(wout8_52),
                    .aout1(aout9_52), .aout2(aout10_52), .aout3(aout11_52), .aout4(aout12_52),
                    .wout1(wout12_49), .wout2(wout12_50), .wout3(wout12_51), .wout4(wout12_52),
                    .sout11(sout9_49), .sout12(sout9_50), .sout13(sout9_51), .sout14(sout9_52),
                    .sout21(sout10_49), .sout22(sout10_50), .sout23(sout10_51), .sout24(sout10_52),
                    .sout31(sout11_49), .sout32(sout11_50), .sout33(sout11_51), .sout34(sout11_52),
                    .sout41(sout12_49), .sout42(sout12_50), .sout43(sout12_51), .sout44(sout12_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_3_14 (.clk(clk), .rst(rst),
                    .ain1(aout9_52), .ain2(aout10_52), .ain3(aout11_52), .ain4(aout12_52),
                    .win1(wout8_53), .win2(wout8_54), .win3(wout8_55), .win4(wout8_56),
                    .aout1(aout9_56), .aout2(aout10_56), .aout3(aout11_56), .aout4(aout12_56),
                    .wout1(wout12_53), .wout2(wout12_54), .wout3(wout12_55), .wout4(wout12_56),
                    .sout11(sout9_53), .sout12(sout9_54), .sout13(sout9_55), .sout14(sout9_56),
                    .sout21(sout10_53), .sout22(sout10_54), .sout23(sout10_55), .sout24(sout10_56),
                    .sout31(sout11_53), .sout32(sout11_54), .sout33(sout11_55), .sout34(sout11_56),
                    .sout41(sout12_53), .sout42(sout12_54), .sout43(sout12_55), .sout44(sout12_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_3_15 (.clk(clk), .rst(rst),
                    .ain1(aout9_56), .ain2(aout10_56), .ain3(aout11_56), .ain4(aout12_56),
                    .win1(wout8_57), .win2(wout8_58), .win3(wout8_59), .win4(wout8_60),
                    .aout1(aout9_60), .aout2(aout10_60), .aout3(aout11_60), .aout4(aout12_60),
                    .wout1(wout12_57), .wout2(wout12_58), .wout3(wout12_59), .wout4(wout12_60),
                    .sout11(sout9_57), .sout12(sout9_58), .sout13(sout9_59), .sout14(sout9_60),
                    .sout21(sout10_57), .sout22(sout10_58), .sout23(sout10_59), .sout24(sout10_60),
                    .sout31(sout11_57), .sout32(sout11_58), .sout33(sout11_59), .sout34(sout11_60),
                    .sout41(sout12_57), .sout42(sout12_58), .sout43(sout12_59), .sout44(sout12_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_3_16 (.clk(clk), .rst(rst),
                    .ain1(aout9_60), .ain2(aout10_60), .ain3(aout11_60), .ain4(aout12_60),
                    .win1(wout8_61), .win2(wout8_62), .win3(wout8_63), .win4(wout8_64),
                    .aout1(aout9_64), .aout2(aout10_64), .aout3(aout11_64), .aout4(aout12_64),
                    .wout1(wout12_61), .wout2(wout12_62), .wout3(wout12_63), .wout4(wout12_64),
                    .sout11(sout9_61), .sout12(sout9_62), .sout13(sout9_63), .sout14(sout9_64),
                    .sout21(sout10_61), .sout22(sout10_62), .sout23(sout10_63), .sout24(sout10_64),
                    .sout31(sout11_61), .sout32(sout11_62), .sout33(sout11_63), .sout34(sout11_64),
                    .sout41(sout12_61), .sout42(sout12_62), .sout43(sout12_63), .sout44(sout12_64)
                    ); //4x4 MAC array
               
                    
                    
    //row4
    mac_array_4x4 mac_array_4x4_41 (.clk(clk), .rst(rst),
                    .ain1(ain13), .ain2(ain14), .ain3(ain15), .ain4(ain16),
                    .win1(wout12_1), .win2(wout12_2), .win3(wout12_3), .win4(wout12_4),
                    .aout1(aout13_4), .aout2(aout14_4), .aout3(aout15_4), .aout4(aout16_4),
                    .wout1(wout16_1), .wout2(wout16_2), .wout3(wout16_3), .wout4(wout16_4),
                    .sout11(sout13_1), .sout12(sout13_2), .sout13(sout13_3), .sout14(sout13_4),
                    .sout21(sout14_1), .sout22(sout14_2), .sout23(sout14_3), .sout24(sout14_4),
                    .sout31(sout15_1), .sout32(sout15_2), .sout33(sout15_3), .sout34(sout15_4),
                    .sout41(sout16_1), .sout42(sout16_2), .sout43(sout16_3), .sout44(sout16_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_42 (.clk(clk), .rst(rst),
                    .ain1(aout13_4), .ain2(aout14_4), .ain3(aout15_4), .ain4(aout16_4),
                    .win1(wout12_5), .win2(wout12_6), .win3(wout12_7), .win4(wout12_8),
                    .aout1(aout13_8), .aout2(aout14_8), .aout3(aout15_8), .aout4(aout16_8),
                    .wout1(wout16_5), .wout2(wout16_6), .wout3(wout16_7), .wout4(wout16_8),
                    .sout11(sout13_5), .sout12(sout13_6), .sout13(sout13_7), .sout14(sout13_8),
                    .sout21(sout14_5), .sout22(sout14_6), .sout23(sout14_7), .sout24(sout14_8),
                    .sout31(sout15_5), .sout32(sout15_6), .sout33(sout15_7), .sout34(sout15_8),
                    .sout41(sout16_5), .sout42(sout16_6), .sout43(sout16_7), .sout44(sout16_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_43 (.clk(clk), .rst(rst),
                    .ain1(aout13_8), .ain2(aout14_8), .ain3(aout15_8), .ain4(aout16_8),
                    .win1(wout12_9), .win2(wout12_10), .win3(wout12_11), .win4(wout12_12),
                    .aout1(aout13_12), .aout2(aout14_12), .aout3(aout15_12), .aout4(aout16_12),
                    .wout1(wout16_9), .wout2(wout16_10), .wout3(wout16_11), .wout4(wout16_12),
                    .sout11(sout13_9), .sout12(sout13_10), .sout13(sout13_11), .sout14(sout13_12),
                    .sout21(sout14_9), .sout22(sout14_10), .sout23(sout14_11), .sout24(sout14_12),
                    .sout31(sout15_9), .sout32(sout15_10), .sout33(sout15_11), .sout34(sout15_12),
                    .sout41(sout16_9), .sout42(sout16_10), .sout43(sout16_11), .sout44(sout16_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_44 (.clk(clk), .rst(rst),
                    .ain1(aout13_12), .ain2(aout14_12), .ain3(aout15_12), .ain4(aout16_12),
                    .win1(wout12_13), .win2(wout12_14), .win3(wout12_15), .win4(wout12_16),
                    .aout1(aout13_16), .aout2(aout14_16), .aout3(aout15_16), .aout4(aout16_16),
                    .wout1(wout16_13), .wout2(wout16_14), .wout3(wout16_15), .wout4(wout16_16),
                    .sout11(sout13_13), .sout12(sout13_14), .sout13(sout13_15), .sout14(sout13_16),
                    .sout21(sout14_13), .sout22(sout14_14), .sout23(sout14_15), .sout24(sout14_16),
                    .sout31(sout15_13), .sout32(sout15_14), .sout33(sout15_15), .sout34(sout15_16),
                    .sout41(sout16_13), .sout42(sout16_14), .sout43(sout16_15), .sout44(sout16_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_45 (.clk(clk), .rst(rst),
                    .ain1(aout13_16), .ain2(aout14_16), .ain3(aout15_16), .ain4(aout16_16),
                    .win1(wout12_17), .win2(wout12_18), .win3(wout12_19), .win4(wout12_20),
                    .aout1(aout13_20), .aout2(aout14_20), .aout3(aout15_20), .aout4(aout16_20),
                    .wout1(wout16_17), .wout2(wout16_18), .wout3(wout16_19), .wout4(wout16_20),
                    .sout11(sout13_17), .sout12(sout13_18), .sout13(sout13_19), .sout14(sout13_20),
                    .sout21(sout14_17), .sout22(sout14_18), .sout23(sout14_19), .sout24(sout14_20),
                    .sout31(sout15_17), .sout32(sout15_18), .sout33(sout15_19), .sout34(sout15_20),
                    .sout41(sout16_17), .sout42(sout16_18), .sout43(sout16_19), .sout44(sout16_20)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_46 (.clk(clk), .rst(rst),
                    .ain1(aout13_20), .ain2(aout14_20), .ain3(aout15_20), .ain4(aout16_20),
                    .win1(wout12_21), .win2(wout12_22), .win3(wout12_23), .win4(wout12_24),
                    .aout1(aout13_24), .aout2(aout14_24), .aout3(aout15_24), .aout4(aout16_24),
                    .wout1(wout16_21), .wout2(wout16_22), .wout3(wout16_23), .wout4(wout16_24),
                    .sout11(sout13_21), .sout12(sout13_22), .sout13(sout13_23), .sout14(sout13_24),
                    .sout21(sout14_21), .sout22(sout14_22), .sout23(sout14_23), .sout24(sout14_24),
                    .sout31(sout15_21), .sout32(sout15_22), .sout33(sout15_23), .sout34(sout15_24),
                    .sout41(sout16_21), .sout42(sout16_22), .sout43(sout16_23), .sout44(sout16_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_47 (.clk(clk), .rst(rst),
                    .ain1(aout13_24), .ain2(aout14_24), .ain3(aout15_24), .ain4(aout16_24),
                    .win1(wout12_25), .win2(wout12_26), .win3(wout12_27), .win4(wout12_28),
                    .aout1(aout13_28), .aout2(aout14_28), .aout3(aout15_28), .aout4(aout16_28),
                    .wout1(wout16_25), .wout2(wout16_26), .wout3(wout16_27), .wout4(wout16_28),
                    .sout11(sout13_25), .sout12(sout13_26), .sout13(sout13_27), .sout14(sout13_28),
                    .sout21(sout14_25), .sout22(sout14_26), .sout23(sout14_27), .sout24(sout14_28),
                    .sout31(sout15_25), .sout32(sout15_26), .sout33(sout15_27), .sout34(sout15_28),
                    .sout41(sout16_25), .sout42(sout16_26), .sout43(sout16_27), .sout44(sout16_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_48 (.clk(clk), .rst(rst),
                    .ain1(aout13_28), .ain2(aout14_28), .ain3(aout15_28), .ain4(aout16_28),
                    .win1(wout12_29), .win2(wout12_30), .win3(wout12_31), .win4(wout12_32),
                    .aout1(aout13_32), .aout2(aout14_32), .aout3(aout15_32), .aout4(aout16_32),
                    .wout1(wout16_29), .wout2(wout16_30), .wout3(wout16_31), .wout4(wout16_32),
                    .sout11(sout13_29), .sout12(sout13_30), .sout13(sout13_31), .sout14(sout13_32),
                    .sout21(sout14_29), .sout22(sout14_30), .sout23(sout14_31), .sout24(sout14_32),
                    .sout31(sout15_29), .sout32(sout15_30), .sout33(sout15_31), .sout34(sout15_32),
                    .sout41(sout16_29), .sout42(sout16_30), .sout43(sout16_31), .sout44(sout16_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_49 (.clk(clk), .rst(rst),
                    .ain1(aout13_32), .ain2(aout14_32), .ain3(aout15_32), .ain4(aout16_32),
                    .win1(wout12_33), .win2(wout12_34), .win3(wout12_35), .win4(wout12_36),
                    .aout1(aout13_36), .aout2(aout14_36), .aout3(aout15_36), .aout4(aout16_36),
                    .wout1(wout16_33), .wout2(wout16_34), .wout3(wout16_35), .wout4(wout16_36),
                    .sout11(sout13_33), .sout12(sout13_34), .sout13(sout13_35), .sout14(sout13_36),
                    .sout21(sout14_33), .sout22(sout14_34), .sout23(sout14_35), .sout24(sout14_36),
                    .sout31(sout15_33), .sout32(sout15_34), .sout33(sout15_35), .sout34(sout15_36),
                    .sout41(sout16_33), .sout42(sout16_34), .sout43(sout16_35), .sout44(sout16_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_4_10 (.clk(clk), .rst(rst),
                    .ain1(aout13_36), .ain2(aout14_36), .ain3(aout15_36), .ain4(aout16_36),
                    .win1(wout12_37), .win2(wout12_38), .win3(wout12_39), .win4(wout12_40),
                    .aout1(aout13_40), .aout2(aout14_40), .aout3(aout15_40), .aout4(aout16_40),
                    .wout1(wout16_37), .wout2(wout16_38), .wout3(wout16_39), .wout4(wout16_40),
                    .sout11(sout13_37), .sout12(sout13_38), .sout13(sout13_39), .sout14(sout13_40),
                    .sout21(sout14_37), .sout22(sout14_38), .sout23(sout14_39), .sout24(sout14_40),
                    .sout31(sout15_37), .sout32(sout15_38), .sout33(sout15_39), .sout34(sout15_40),
                    .sout41(sout16_37), .sout42(sout16_38), .sout43(sout16_39), .sout44(sout16_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_4_11 (.clk(clk), .rst(rst),
                    .ain1(aout13_40), .ain2(aout14_40), .ain3(aout15_40), .ain4(aout16_40),
                    .win1(wout12_41), .win2(wout12_42), .win3(wout12_43), .win4(wout12_44),
                    .aout1(aout13_44), .aout2(aout14_44), .aout3(aout15_44), .aout4(aout16_44),
                    .wout1(wout16_41), .wout2(wout16_42), .wout3(wout16_43), .wout4(wout16_44),
                    .sout11(sout13_41), .sout12(sout13_42), .sout13(sout13_43), .sout14(sout13_44),
                    .sout21(sout14_41), .sout22(sout14_42), .sout23(sout14_43), .sout24(sout14_44),
                    .sout31(sout15_41), .sout32(sout15_42), .sout33(sout15_43), .sout34(sout15_44),
                    .sout41(sout16_41), .sout42(sout16_42), .sout43(sout16_43), .sout44(sout16_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_4_12 (.clk(clk), .rst(rst),
                    .ain1(aout13_44), .ain2(aout14_44), .ain3(aout15_44), .ain4(aout16_44),
                    .win1(wout12_45), .win2(wout12_46), .win3(wout12_47), .win4(wout12_48),
                    .aout1(aout13_48), .aout2(aout14_48), .aout3(aout15_48), .aout4(aout16_48),
                    .wout1(wout16_45), .wout2(wout16_46), .wout3(wout16_47), .wout4(wout16_48),
                    .sout11(sout13_45), .sout12(sout13_46), .sout13(sout13_47), .sout14(sout13_48),
                    .sout21(sout14_45), .sout22(sout14_46), .sout23(sout14_47), .sout24(sout14_48),
                    .sout31(sout15_45), .sout32(sout15_46), .sout33(sout15_47), .sout34(sout15_48),
                    .sout41(sout16_45), .sout42(sout16_46), .sout43(sout16_47), .sout44(sout16_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_4_13 (.clk(clk), .rst(rst),
                    .ain1(aout13_48), .ain2(aout14_48), .ain3(aout15_48), .ain4(aout16_48),
                    .win1(wout12_49), .win2(wout12_50), .win3(wout12_51), .win4(wout12_52),
                    .aout1(aout13_52), .aout2(aout14_52), .aout3(aout15_52), .aout4(aout16_52),
                    .wout1(wout16_49), .wout2(wout16_50), .wout3(wout16_51), .wout4(wout16_52),
                    .sout11(sout13_49), .sout12(sout13_50), .sout13(sout13_51), .sout14(sout13_52),
                    .sout21(sout14_49), .sout22(sout14_50), .sout23(sout14_51), .sout24(sout14_52),
                    .sout31(sout15_49), .sout32(sout15_50), .sout33(sout15_51), .sout34(sout15_52),
                    .sout41(sout16_49), .sout42(sout16_50), .sout43(sout16_51), .sout44(sout16_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_4_14 (.clk(clk), .rst(rst),
                    .ain1(aout13_52), .ain2(aout14_52), .ain3(aout15_52), .ain4(aout16_52),
                    .win1(wout12_53), .win2(wout12_54), .win3(wout12_55), .win4(wout12_56),
                    .aout1(aout13_56), .aout2(aout14_56), .aout3(aout15_56), .aout4(aout16_56),
                    .wout1(wout16_53), .wout2(wout16_54), .wout3(wout16_55), .wout4(wout16_56),
                    .sout11(sout13_53), .sout12(sout13_54), .sout13(sout13_55), .sout14(sout13_56),
                    .sout21(sout14_53), .sout22(sout14_54), .sout23(sout14_55), .sout24(sout14_56),
                    .sout31(sout15_53), .sout32(sout15_54), .sout33(sout15_55), .sout34(sout15_56),
                    .sout41(sout16_53), .sout42(sout16_54), .sout43(sout16_55), .sout44(sout16_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_4_15 (.clk(clk), .rst(rst),
                    .ain1(aout13_56), .ain2(aout14_56), .ain3(aout15_56), .ain4(aout16_56),
                    .win1(wout12_57), .win2(wout12_58), .win3(wout12_59), .win4(wout12_60),
                    .aout1(aout13_60), .aout2(aout14_60), .aout3(aout15_60), .aout4(aout16_60),
                    .wout1(wout16_57), .wout2(wout16_58), .wout3(wout16_59), .wout4(wout16_60),
                    .sout11(sout13_57), .sout12(sout13_58), .sout13(sout13_59), .sout14(sout13_60),
                    .sout21(sout14_57), .sout22(sout14_58), .sout23(sout14_59), .sout24(sout14_60),
                    .sout31(sout15_57), .sout32(sout15_58), .sout33(sout15_59), .sout34(sout15_60),
                    .sout41(sout16_57), .sout42(sout16_58), .sout43(sout16_59), .sout44(sout16_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_4_16 (.clk(clk), .rst(rst),
                    .ain1(aout13_60), .ain2(aout14_60), .ain3(aout15_60), .ain4(aout16_60),
                    .win1(wout12_61), .win2(wout12_62), .win3(wout12_63), .win4(wout12_64),
                    .aout1(aout13_64), .aout2(aout14_64), .aout3(aout15_64), .aout4(aout16_64),
                    .wout1(wout16_61), .wout2(wout16_62), .wout3(wout16_63), .wout4(wout16_64),
                    .sout11(sout13_61), .sout12(sout13_62), .sout13(sout13_63), .sout14(sout13_64),
                    .sout21(sout14_61), .sout22(sout14_62), .sout23(sout14_63), .sout24(sout14_64),
                    .sout31(sout15_61), .sout32(sout15_62), .sout33(sout15_63), .sout34(sout15_64),
                    .sout41(sout16_61), .sout42(sout16_62), .sout43(sout16_63), .sout44(sout16_64)
                    ); //4x4 MAC array
                    
    
    //row5
    mac_array_4x4 mac_array_4x4_51 (.clk(clk), .rst(rst),
                    .ain1(ain17), .ain2(ain18), .ain3(ain19), .ain4(ain20),
                    .win1(wout16_1), .win2(wout16_2), .win3(wout16_3), .win4(wout16_4),
                    .aout1(aout17_4), .aout2(aout18_4), .aout3(aout19_4), .aout4(aout20_4),
                    .wout1(wout20_1), .wout2(wout20_2), .wout3(wout20_3), .wout4(wout20_4),
                    .sout11(sout17_1), .sout12(sout17_2), .sout13(sout17_3), .sout14(sout17_4),
                    .sout21(sout18_1), .sout22(sout18_2), .sout23(sout18_3), .sout24(sout18_4),
                    .sout31(sout19_1), .sout32(sout19_2), .sout33(sout19_3), .sout34(sout19_4),
                    .sout41(sout20_1), .sout42(sout20_2), .sout43(sout20_3), .sout44(sout20_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_52 (.clk(clk), .rst(rst),
                    .ain1(aout17_4), .ain2(aout18_4), .ain3(aout18_4), .ain4(aout20_4),
                    .win1(wout16_5), .win2(wout16_6), .win3(wout16_7), .win4(wout16_8),
                    .aout1(aout17_8), .aout2(aout18_8), .aout3(aout19_8), .aout4(aout20_8),
                    .wout1(wout20_5), .wout2(wout20_6), .wout3(wout20_7), .wout4(wout20_8),
                    .sout11(sout17_5), .sout12(sout17_6), .sout13(sout17_7), .sout14(sout17_8),
                    .sout21(sout18_5), .sout22(sout18_6), .sout23(sout18_7), .sout24(sout18_8),
                    .sout31(sout19_5), .sout32(sout19_6), .sout33(sout19_7), .sout34(sout19_8),
                    .sout41(sout20_5), .sout42(sout20_6), .sout43(sout20_7), .sout44(sout20_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_53 (.clk(clk), .rst(rst),
                    .ain1(aout17_8), .ain2(aout18_8), .ain3(aout19_8), .ain4(aout20_8),
                    .win1(wout16_9), .win2(wout16_10), .win3(wout16_11), .win4(wout16_12),
                    .aout1(aout17_12), .aout2(aout18_12), .aout3(aout19_12), .aout4(aout20_12),
                    .wout1(wout20_9), .wout2(wout20_10), .wout3(wout20_11), .wout4(wout20_12),
                    .sout11(sout17_9), .sout12(sout17_10), .sout13(sout17_11), .sout14(sout17_12),
                    .sout21(sout18_9), .sout22(sout18_10), .sout23(sout18_11), .sout24(sout18_12),
                    .sout31(sout19_9), .sout32(sout19_10), .sout33(sout19_11), .sout34(sout19_12),
                    .sout41(sout20_9), .sout42(sout20_10), .sout43(sout20_11), .sout44(sout20_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_54 (.clk(clk), .rst(rst),
                    .ain1(aout17_12), .ain2(aout18_12), .ain3(aout19_12), .ain4(aout20_12),
                    .win1(wout16_13), .win2(wout16_14), .win3(wout16_15), .win4(wout16_16),
                    .aout1(aout17_16), .aout2(aout18_16), .aout3(aout19_16), .aout4(aout20_16),
                    .wout1(wout20_13), .wout2(wout20_14), .wout3(wout20_15), .wout4(wout20_16),
                    .sout11(sout17_13), .sout12(sout17_14), .sout13(sout17_15), .sout14(sout17_16),
                    .sout21(sout18_13), .sout22(sout18_14), .sout23(sout18_15), .sout24(sout18_16),
                    .sout31(sout19_13), .sout32(sout19_14), .sout33(sout19_15), .sout34(sout19_16),
                    .sout41(sout20_13), .sout42(sout20_14), .sout43(sout20_15), .sout44(sout20_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_55 (.clk(clk), .rst(rst),
                    .ain1(aout17_16), .ain2(aout18_16), .ain3(aout19_16), .ain4(aout20_16),
                    .win1(wout16_17), .win2(wout16_18), .win3(wout16_19), .win4(wout16_20),
                    .aout1(aout17_20), .aout2(aout18_20), .aout3(aout19_20), .aout4(aout20_20),
                    .wout1(wout20_17), .wout2(wout20_18), .wout3(wout20_19), .wout4(wout20_20),
                    .sout11(sout17_17), .sout12(sout17_18), .sout13(sout17_19), .sout14(sout17_20),
                    .sout21(sout18_17), .sout22(sout18_18), .sout23(sout18_19), .sout24(sout18_20),
                    .sout31(sout19_17), .sout32(sout19_18), .sout33(sout19_19), .sout34(sout19_20),
                    .sout41(sout20_17), .sout42(sout20_18), .sout43(sout20_19), .sout44(sout20_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_56 (.clk(clk), .rst(rst),
                    .ain1(aout17_20), .ain2(aout18_20), .ain3(aout19_20), .ain4(aout20_20),
                    .win1(wout16_21), .win2(wout16_22), .win3(wout16_23), .win4(wout16_24),
                    .aout1(aout17_24), .aout2(aout18_24), .aout3(aout19_24), .aout4(aout20_24),
                    .wout1(wout20_21), .wout2(wout20_22), .wout3(wout20_23), .wout4(wout20_24),
                    .sout11(sout17_21), .sout12(sout17_22), .sout13(sout17_23), .sout14(sout17_24),
                    .sout21(sout18_21), .sout22(sout18_22), .sout23(sout18_23), .sout24(sout18_24),
                    .sout31(sout19_21), .sout32(sout19_22), .sout33(sout19_23), .sout34(sout19_24),
                    .sout41(sout20_21), .sout42(sout20_22), .sout43(sout20_23), .sout44(sout20_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_57 (.clk(clk), .rst(rst),
                    .ain1(aout17_24), .ain2(aout18_24), .ain3(aout19_24), .ain4(aout20_24),
                    .win1(wout16_25), .win2(wout16_26), .win3(wout16_27), .win4(wout16_28),
                    .aout1(aout17_28), .aout2(aout18_28), .aout3(aout19_28), .aout4(aout20_28),
                    .wout1(wout20_25), .wout2(wout20_26), .wout3(wout20_27), .wout4(wout20_28),
                    .sout11(sout17_25), .sout12(sout17_26), .sout13(sout17_27), .sout14(sout17_28),
                    .sout21(sout18_25), .sout22(sout18_26), .sout23(sout18_27), .sout24(sout18_28),
                    .sout31(sout19_25), .sout32(sout19_26), .sout33(sout19_27), .sout34(sout19_28),
                    .sout41(sout20_25), .sout42(sout20_26), .sout43(sout20_27), .sout44(sout20_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_58 (.clk(clk), .rst(rst),
                    .ain1(aout17_28), .ain2(aout18_28), .ain3(aout19_28), .ain4(aout20_28),
                    .win1(wout16_29), .win2(wout16_30), .win3(wout16_31), .win4(wout16_32),
                    .aout1(aout17_32), .aout2(aout18_32), .aout3(aout19_32), .aout4(aout20_32),
                    .wout1(wout20_29), .wout2(wout20_30), .wout3(wout20_31), .wout4(wout20_32),
                    .sout11(sout17_29), .sout12(sout17_30), .sout13(sout17_31), .sout14(sout17_32),
                    .sout21(sout18_29), .sout22(sout18_30), .sout23(sout18_31), .sout24(sout18_32),
                    .sout31(sout19_29), .sout32(sout19_30), .sout33(sout19_31), .sout34(sout19_32),
                    .sout41(sout20_29), .sout42(sout20_30), .sout43(sout20_31), .sout44(sout20_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_59 (.clk(clk), .rst(rst),
                    .ain1(aout17_32), .ain2(aout18_32), .ain3(aout19_32), .ain4(aout20_32),
                    .win1(wout16_33), .win2(wout16_34), .win3(wout16_35), .win4(wout16_36),
                    .aout1(aout17_36), .aout2(aout18_36), .aout3(aout19_36), .aout4(aout20_36),
                    .wout1(wout20_33), .wout2(wout20_34), .wout3(wout20_35), .wout4(wout20_36),
                    .sout11(sout17_33), .sout12(sout17_34), .sout13(sout17_35), .sout14(sout17_36),
                    .sout21(sout18_33), .sout22(sout18_34), .sout23(sout18_35), .sout24(sout18_36),
                    .sout31(sout19_33), .sout32(sout19_34), .sout33(sout19_35), .sout34(sout19_36),
                    .sout41(sout20_33), .sout42(sout20_34), .sout43(sout20_35), .sout44(sout20_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_5_10 (.clk(clk), .rst(rst),
                    .ain1(aout17_36), .ain2(aout18_36), .ain3(aout19_36), .ain4(aout20_36),
                    .win1(wout16_37), .win2(wout16_38), .win3(wout16_39), .win4(wout16_40),
                    .aout1(aout17_40), .aout2(aout18_40), .aout3(aout19_40), .aout4(aout20_40),
                    .wout1(wout20_37), .wout2(wout20_38), .wout3(wout20_39), .wout4(wout20_40),
                    .sout11(sout17_37), .sout12(sout17_38), .sout13(sout17_39), .sout14(sout17_40),
                    .sout21(sout18_37), .sout22(sout18_38), .sout23(sout18_39), .sout24(sout18_40),
                    .sout31(sout19_37), .sout32(sout19_38), .sout33(sout19_39), .sout34(sout19_40),
                    .sout41(sout20_37), .sout42(sout20_38), .sout43(sout20_39), .sout44(sout20_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_5_11 (.clk(clk), .rst(rst),
                    .ain1(aout17_40), .ain2(aout18_40), .ain3(aout19_40), .ain4(aout20_40),
                    .win1(wout16_41), .win2(wout16_42), .win3(wout16_43), .win4(wout16_44),
                    .aout1(aout17_44), .aout2(aout18_44), .aout3(aout19_44), .aout4(aout20_44),
                    .wout1(wout20_41), .wout2(wout20_42), .wout3(wout20_43), .wout4(wout20_44),
                    .sout11(sout17_41), .sout12(sout17_42), .sout13(sout17_43), .sout14(sout17_44),
                    .sout21(sout18_41), .sout22(sout18_42), .sout23(sout18_43), .sout24(sout18_44),
                    .sout31(sout19_41), .sout32(sout19_42), .sout33(sout19_43), .sout34(sout19_44),
                    .sout41(sout20_41), .sout42(sout20_42), .sout43(sout20_43), .sout44(sout20_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_5_12 (.clk(clk), .rst(rst),
                    .ain1(aout17_44), .ain2(aout18_44), .ain3(aout19_44), .ain4(aout20_44),
                    .win1(wout16_45), .win2(wout16_46), .win3(wout16_47), .win4(wout16_48),
                    .aout1(aout17_48), .aout2(aout18_48), .aout3(aout19_48), .aout4(aout20_48),
                    .wout1(wout20_45), .wout2(wout20_46), .wout3(wout20_47), .wout4(wout20_48),
                    .sout11(sout17_45), .sout12(sout17_46), .sout13(sout17_47), .sout14(sout17_48),
                    .sout21(sout18_45), .sout22(sout18_46), .sout23(sout18_47), .sout24(sout18_48),
                    .sout31(sout19_45), .sout32(sout19_46), .sout33(sout19_47), .sout34(sout19_48),
                    .sout41(sout20_45), .sout42(sout20_46), .sout43(sout20_47), .sout44(sout20_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_5_13 (.clk(clk), .rst(rst),
                    .ain1(aout17_48), .ain2(aout18_48), .ain3(aout19_48), .ain4(aout20_48),
                    .win1(wout16_49), .win2(wout16_50), .win3(wout16_51), .win4(wout16_52),
                    .aout1(aout17_52), .aout2(aout18_52), .aout3(aout19_52), .aout4(aout20_52),
                    .wout1(wout20_49), .wout2(wout20_50), .wout3(wout20_51), .wout4(wout20_52),
                    .sout11(sout17_49), .sout12(sout17_50), .sout13(sout17_51), .sout14(sout17_52),
                    .sout21(sout18_49), .sout22(sout18_50), .sout23(sout18_51), .sout24(sout18_52),
                    .sout31(sout19_49), .sout32(sout19_50), .sout33(sout19_51), .sout34(sout19_52),
                    .sout41(sout20_49), .sout42(sout20_50), .sout43(sout20_51), .sout44(sout20_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_5_14 (.clk(clk), .rst(rst),
                    .ain1(aout17_52), .ain2(aout18_52), .ain3(aout19_52), .ain4(aout20_52),
                    .win1(wout16_53), .win2(wout16_54), .win3(wout16_55), .win4(wout16_56),
                    .aout1(aout17_56), .aout2(aout18_56), .aout3(aout19_56), .aout4(aout20_56),
                    .wout1(wout20_53), .wout2(wout20_54), .wout3(wout20_55), .wout4(wout20_56),
                    .sout11(sout17_53), .sout12(sout17_54), .sout13(sout17_55), .sout14(sout17_56),
                    .sout21(sout18_53), .sout22(sout18_54), .sout23(sout18_55), .sout24(sout18_56),
                    .sout31(sout19_53), .sout32(sout19_54), .sout33(sout19_55), .sout34(sout19_56),
                    .sout41(sout20_53), .sout42(sout20_54), .sout43(sout20_55), .sout44(sout20_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_5_15 (.clk(clk), .rst(rst),
                    .ain1(aout17_56), .ain2(aout18_56), .ain3(aout19_56), .ain4(aout20_56),
                    .win1(wout16_57), .win2(wout16_58), .win3(wout16_59), .win4(wout16_60),
                    .aout1(aout17_60), .aout2(aout18_60), .aout3(aout19_60), .aout4(aout20_60),
                    .wout1(wout20_57), .wout2(wout20_58), .wout3(wout20_59), .wout4(wout20_60),
                    .sout11(sout17_57), .sout12(sout17_58), .sout13(sout17_59), .sout14(sout17_60),
                    .sout21(sout18_57), .sout22(sout18_58), .sout23(sout18_59), .sout24(sout18_60),
                    .sout31(sout19_57), .sout32(sout19_58), .sout33(sout19_59), .sout34(sout19_60),
                    .sout41(sout20_57), .sout42(sout20_58), .sout43(sout20_59), .sout44(sout20_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_5_16 (.clk(clk), .rst(rst),
                    .ain1(aout17_60), .ain2(aout18_60), .ain3(aout19_60), .ain4(aout20_60),
                    .win1(wout16_61), .win2(wout16_62), .win3(wout16_63), .win4(wout16_64),
                    .aout1(aout17_64), .aout2(aout18_64), .aout3(aout19_64), .aout4(aout20_64),
                    .wout1(wout20_61), .wout2(wout20_62), .wout3(wout20_63), .wout4(wout20_64),
                    .sout11(sout17_61), .sout12(sout17_62), .sout13(sout17_63), .sout14(sout17_64),
                    .sout21(sout18_61), .sout22(sout18_62), .sout23(sout18_63), .sout24(sout18_64),
                    .sout31(sout19_61), .sout32(sout19_62), .sout33(sout19_63), .sout34(sout19_64),
                    .sout41(sout20_61), .sout42(sout20_62), .sout43(sout20_63), .sout44(sout20_64)
                    ); //4x4 MAC array
    
    
    //row6
    mac_array_4x4 mac_array_4x4_61 (.clk(clk), .rst(rst),
                    .ain1(ain21), .ain2(ain22), .ain3(ain23), .ain4(ain24),
                    .win1(wout20_1), .win2(wout20_2), .win3(wout20_3), .win4(wout20_4),
                    .aout1(aout21_4), .aout2(aout22_4), .aout3(aout23_4), .aout4(aout24_4),
                    .wout1(wout24_1), .wout2(wout24_2), .wout3(wout24_3), .wout4(wout24_4),
                    .sout11(sout21_1), .sout12(sout21_2), .sout13(sout21_3), .sout14(sout21_4),
                    .sout21(sout22_1), .sout22(sout22_2), .sout23(sout22_3), .sout24(sout22_4),
                    .sout31(sout23_1), .sout32(sout23_2), .sout33(sout23_3), .sout34(sout23_4),
                    .sout41(sout24_1), .sout42(sout24_2), .sout43(sout24_3), .sout44(sout24_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_62 (.clk(clk), .rst(rst),
                    .ain1(aout21_4), .ain2(aout22_4), .ain3(aout23_4), .ain4(aout24_4),
                    .win1(wout20_5), .win2(wout20_6), .win3(wout20_7), .win4(wout20_8),
                    .aout1(aout21_8), .aout2(aout22_8), .aout3(aout23_8), .aout4(aout24_8),
                    .wout1(wout24_5), .wout2(wout24_6), .wout3(wout24_7), .wout4(wout24_8),
                    .sout11(sout21_5), .sout12(sout21_6), .sout13(sout21_7), .sout14(sout21_8),
                    .sout21(sout22_5), .sout22(sout22_6), .sout23(sout22_7), .sout24(sout22_8),
                    .sout31(sout23_5), .sout32(sout23_6), .sout33(sout23_7), .sout34(sout23_8),
                    .sout41(sout24_5), .sout42(sout24_6), .sout43(sout24_7), .sout44(sout24_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_63 (.clk(clk), .rst(rst),
                    .ain1(aout21_8), .ain2(aout22_8), .ain3(aout23_8), .ain4(aout24_8),
                    .win1(wout20_9), .win2(wout20_10), .win3(wout20_11), .win4(wout20_12),
                    .aout1(aout21_12), .aout2(aout22_12), .aout3(aout23_12), .aout4(aout24_12),
                    .wout1(wout24_9), .wout2(wout24_10), .wout3(wout24_11), .wout4(wout24_12),
                    .sout11(sout21_9), .sout12(sout21_10), .sout13(sout21_11), .sout14(sout21_12),
                    .sout21(sout22_9), .sout22(sout22_10), .sout23(sout22_11), .sout24(sout22_12),
                    .sout31(sout23_9), .sout32(sout23_10), .sout33(sout23_11), .sout34(sout23_12),
                    .sout41(sout24_9), .sout42(sout24_10), .sout43(sout24_11), .sout44(sout24_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_64 (.clk(clk), .rst(rst),
                    .ain1(aout21_12), .ain2(aout22_12), .ain3(aout23_12), .ain4(aout24_12),
                    .win1(wout20_13), .win2(wout20_14), .win3(wout20_15), .win4(wout20_16),
                    .aout1(aout21_16), .aout2(aout22_16), .aout3(aout23_16), .aout4(aout24_16),
                    .wout1(wout24_13), .wout2(wout24_14), .wout3(wout24_15), .wout4(wout24_16),
                    .sout11(sout21_13), .sout12(sout21_14), .sout13(sout21_15), .sout14(sout21_16),
                    .sout21(sout22_13), .sout22(sout22_14), .sout23(sout22_15), .sout24(sout22_16),
                    .sout31(sout23_13), .sout32(sout23_14), .sout33(sout23_15), .sout34(sout23_16),
                    .sout41(sout24_13), .sout42(sout24_14), .sout43(sout24_15), .sout44(sout24_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_65 (.clk(clk), .rst(rst),
                    .ain1(aout21_16), .ain2(aout22_16), .ain3(aout23_16), .ain4(aout24_16),
                    .win1(wout20_17), .win2(wout20_18), .win3(wout20_19), .win4(wout20_20),
                    .aout1(aout21_20), .aout2(aout22_20), .aout3(aout23_20), .aout4(aout24_20),
                    .wout1(wout24_17), .wout2(wout24_18), .wout3(wout24_19), .wout4(wout24_20),
                    .sout11(sout21_17), .sout12(sout21_18), .sout13(sout21_19), .sout14(sout21_20),
                    .sout21(sout22_17), .sout22(sout22_18), .sout23(sout22_19), .sout24(sout22_20),
                    .sout31(sout23_17), .sout32(sout23_18), .sout33(sout23_19), .sout34(sout23_20),
                    .sout41(sout24_17), .sout42(sout24_18), .sout43(sout24_19), .sout44(sout24_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_66 (.clk(clk), .rst(rst),
                    .ain1(aout21_20), .ain2(aout22_20), .ain3(aout23_20), .ain4(aout24_20),
                    .win1(wout20_21), .win2(wout20_22), .win3(wout20_23), .win4(wout20_24),
                    .aout1(aout21_24), .aout2(aout22_24), .aout3(aout23_24), .aout4(aout24_24),
                    .wout1(wout24_21), .wout2(wout24_22), .wout3(wout24_23), .wout4(wout24_24),
                    .sout11(sout21_21), .sout12(sout21_22), .sout13(sout21_23), .sout14(sout21_24),
                    .sout21(sout22_21), .sout22(sout22_22), .sout23(sout22_23), .sout24(sout22_24),
                    .sout31(sout23_21), .sout32(sout23_22), .sout33(sout23_23), .sout34(sout23_24),
                    .sout41(sout24_21), .sout42(sout24_22), .sout43(sout24_23), .sout44(sout24_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_67 (.clk(clk), .rst(rst),
                    .ain1(aout21_24), .ain2(aout22_24), .ain3(aout23_24), .ain4(aout24_24),
                    .win1(wout20_25), .win2(wout20_26), .win3(wout20_27), .win4(wout20_28),
                    .aout1(aout21_28), .aout2(aout22_28), .aout3(aout23_28), .aout4(aout24_28),
                    .wout1(wout24_25), .wout2(wout24_26), .wout3(wout24_27), .wout4(wout24_28),
                    .sout11(sout21_25), .sout12(sout21_26), .sout13(sout21_27), .sout14(sout21_28),
                    .sout21(sout22_25), .sout22(sout22_26), .sout23(sout22_27), .sout24(sout22_28),
                    .sout31(sout23_25), .sout32(sout23_26), .sout33(sout23_27), .sout34(sout23_28),
                    .sout41(sout24_25), .sout42(sout24_26), .sout43(sout24_27), .sout44(sout24_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_68 (.clk(clk), .rst(rst),
                    .ain1(aout21_28), .ain2(aout22_28), .ain3(aout23_28), .ain4(aout24_28),
                    .win1(wout20_29), .win2(wout20_30), .win3(wout20_31), .win4(wout20_32),
                    .aout1(aout21_32), .aout2(aout22_32), .aout3(aout23_32), .aout4(aout24_32),
                    .wout1(wout24_29), .wout2(wout24_30), .wout3(wout24_31), .wout4(wout24_32),
                    .sout11(sout21_29), .sout12(sout21_30), .sout13(sout21_31), .sout14(sout21_32),
                    .sout21(sout22_29), .sout22(sout22_30), .sout23(sout22_31), .sout24(sout22_32),
                    .sout31(sout23_29), .sout32(sout23_30), .sout33(sout23_31), .sout34(sout23_32),
                    .sout41(sout24_29), .sout42(sout24_30), .sout43(sout24_31), .sout44(sout24_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_69 (.clk(clk), .rst(rst),
                    .ain1(aout21_32), .ain2(aout22_32), .ain3(aout23_32), .ain4(aout24_32),
                    .win1(wout20_33), .win2(wout20_34), .win3(wout20_35), .win4(wout20_36),
                    .aout1(aout21_36), .aout2(aout22_36), .aout3(aout23_36), .aout4(aout24_36),
                    .wout1(wout24_33), .wout2(wout24_34), .wout3(wout24_35), .wout4(wout24_36),
                    .sout11(sout21_33), .sout12(sout21_34), .sout13(sout21_35), .sout14(sout21_36),
                    .sout21(sout22_33), .sout22(sout22_34), .sout23(sout22_35), .sout24(sout22_36),
                    .sout31(sout23_33), .sout32(sout23_34), .sout33(sout23_35), .sout34(sout23_36),
                    .sout41(sout24_33), .sout42(sout24_34), .sout43(sout24_35), .sout44(sout24_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_6_10 (.clk(clk), .rst(rst),
                    .ain1(aout21_36), .ain2(aout22_36), .ain3(aout23_36), .ain4(aout24_36),
                    .win1(wout20_37), .win2(wout20_38), .win3(wout20_39), .win4(wout20_40),
                    .aout1(aout21_40), .aout2(aout22_40), .aout3(aout23_40), .aout4(aout24_40),
                    .wout1(wout24_37), .wout2(wout24_38), .wout3(wout24_39), .wout4(wout24_40),
                    .sout11(sout21_37), .sout12(sout21_38), .sout13(sout21_39), .sout14(sout21_40),
                    .sout21(sout22_37), .sout22(sout22_38), .sout23(sout22_39), .sout24(sout22_40),
                    .sout31(sout23_37), .sout32(sout23_38), .sout33(sout23_39), .sout34(sout23_40),
                    .sout41(sout24_37), .sout42(sout24_38), .sout43(sout24_39), .sout44(sout24_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_6_11 (.clk(clk), .rst(rst),
                    .ain1(aout21_40), .ain2(aout22_40), .ain3(aout23_40), .ain4(aout24_40),
                    .win1(wout20_41), .win2(wout20_42), .win3(wout20_43), .win4(wout20_44),
                    .aout1(aout21_44), .aout2(aout22_44), .aout3(aout23_44), .aout4(aout24_44),
                    .wout1(wout24_41), .wout2(wout24_42), .wout3(wout24_43), .wout4(wout24_44),
                    .sout11(sout21_41), .sout12(sout21_42), .sout13(sout21_43), .sout14(sout21_44),
                    .sout21(sout22_41), .sout22(sout22_42), .sout23(sout22_43), .sout24(sout22_44),
                    .sout31(sout23_41), .sout32(sout23_42), .sout33(sout23_43), .sout34(sout23_44),
                    .sout41(sout24_41), .sout42(sout24_42), .sout43(sout24_43), .sout44(sout24_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_6_12 (.clk(clk), .rst(rst),
                    .ain1(aout21_44), .ain2(aout22_44), .ain3(aout23_44), .ain4(aout24_44),
                    .win1(wout20_45), .win2(wout20_46), .win3(wout20_47), .win4(wout20_48),
                    .aout1(aout21_48), .aout2(aout22_48), .aout3(aout23_48), .aout4(aout24_48),
                    .wout1(wout24_45), .wout2(wout24_46), .wout3(wout24_47), .wout4(wout24_48),
                    .sout11(sout21_45), .sout12(sout21_46), .sout13(sout21_47), .sout14(sout21_48),
                    .sout21(sout22_45), .sout22(sout22_46), .sout23(sout22_47), .sout24(sout22_48),
                    .sout31(sout23_45), .sout32(sout23_46), .sout33(sout23_47), .sout34(sout23_48),
                    .sout41(sout24_45), .sout42(sout24_46), .sout43(sout24_47), .sout44(sout24_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_6_13 (.clk(clk), .rst(rst),
                    .ain1(aout21_48), .ain2(aout22_48), .ain3(aout23_48), .ain4(aout24_48),
                    .win1(wout20_49), .win2(wout20_50), .win3(wout20_51), .win4(wout20_52),
                    .aout1(aout21_52), .aout2(aout22_52), .aout3(aout23_52), .aout4(aout24_52),
                    .wout1(wout24_49), .wout2(wout24_50), .wout3(wout24_51), .wout4(wout24_52),
                    .sout11(sout21_49), .sout12(sout21_50), .sout13(sout21_51), .sout14(sout21_52),
                    .sout21(sout22_49), .sout22(sout22_50), .sout23(sout22_51), .sout24(sout22_52),
                    .sout31(sout23_49), .sout32(sout23_50), .sout33(sout23_51), .sout34(sout23_52),
                    .sout41(sout24_49), .sout42(sout24_50), .sout43(sout24_51), .sout44(sout24_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_6_14 (.clk(clk), .rst(rst),
                    .ain1(aout21_52), .ain2(aout22_52), .ain3(aout23_52), .ain4(aout24_52),
                    .win1(wout20_53), .win2(wout20_54), .win3(wout20_55), .win4(wout20_56),
                    .aout1(aout21_56), .aout2(aout22_56), .aout3(aout23_56), .aout4(aout24_56),
                    .wout1(wout24_53), .wout2(wout24_54), .wout3(wout24_55), .wout4(wout24_56),
                    .sout11(sout21_53), .sout12(sout21_54), .sout13(sout21_55), .sout14(sout21_56),
                    .sout21(sout22_53), .sout22(sout22_54), .sout23(sout22_55), .sout24(sout22_56),
                    .sout31(sout23_53), .sout32(sout23_54), .sout33(sout23_55), .sout34(sout23_56),
                    .sout41(sout24_53), .sout42(sout24_54), .sout43(sout24_55), .sout44(sout24_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_6_15 (.clk(clk), .rst(rst),
                    .ain1(aout21_56), .ain2(aout22_56), .ain3(aout23_56), .ain4(aout24_56),
                    .win1(wout20_57), .win2(wout20_58), .win3(wout20_59), .win4(wout20_60),
                    .aout1(aout21_60), .aout2(aout22_60), .aout3(aout23_60), .aout4(aout24_60),
                    .wout1(wout24_57), .wout2(wout24_58), .wout3(wout24_59), .wout4(wout24_60),
                    .sout11(sout17_57), .sout12(sout17_58), .sout13(sout17_59), .sout14(sout17_60),
                    .sout21(sout18_57), .sout22(sout18_58), .sout23(sout18_59), .sout24(sout18_60),
                    .sout31(sout19_57), .sout32(sout19_58), .sout33(sout19_59), .sout34(sout19_60),
                    .sout41(sout20_57), .sout42(sout20_58), .sout43(sout20_59), .sout44(sout20_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_6_16 (.clk(clk), .rst(rst),
                    .ain1(aout21_60), .ain2(aout22_60), .ain3(aout23_60), .ain4(aout24_60),
                    .win1(wout20_61), .win2(wout20_62), .win3(wout20_63), .win4(wout20_64),
                    .aout1(aout21_64), .aout2(aout22_64), .aout3(aout23_64), .aout4(aout24_64),
                    .wout1(wout24_61), .wout2(wout24_62), .wout3(wout24_63), .wout4(wout24_64),
                    .sout11(sout21_61), .sout12(sout21_62), .sout13(sout21_63), .sout14(sout21_64),
                    .sout21(sout22_61), .sout22(sout22_62), .sout23(sout22_63), .sout24(sout22_64),
                    .sout31(sout23_61), .sout32(sout23_62), .sout33(sout23_63), .sout34(sout23_64),
                    .sout41(sout24_61), .sout42(sout24_62), .sout43(sout24_63), .sout44(sout24_64)
                    ); //4x4 MAC array


    //row7
    mac_array_4x4 mac_array_4x4_71 (.clk(clk), .rst(rst),
                    .ain1(ain25), .ain2(ain26), .ain3(ain27), .ain4(ain28),
                    .win1(wout24_1), .win2(wout24_2), .win3(wout24_3), .win4(wout24_4),
                    .aout1(aout25_4), .aout2(aout26_4), .aout3(aout27_4), .aout4(aout28_4),
                    .wout1(wout28_1), .wout2(wout28_2), .wout3(wout28_3), .wout4(wout28_4),
                    .sout11(sout25_1), .sout12(sout25_2), .sout13(sout25_3), .sout14(sout25_4),
                    .sout21(sout26_1), .sout22(sout26_2), .sout23(sout26_3), .sout24(sout26_4),
                    .sout31(sout27_1), .sout32(sout27_2), .sout33(sout27_3), .sout34(sout27_4),
                    .sout41(sout28_1), .sout42(sout28_2), .sout43(sout28_3), .sout44(sout28_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_72 (.clk(clk), .rst(rst),
                    .ain1(aout25_4), .ain2(aout26_4), .ain3(aout27_4), .ain4(aout28_4),
                    .win1(wout24_5), .win2(wout24_6), .win3(wout24_7), .win4(wout24_8),
                    .aout1(aout25_8), .aout2(aout26_8), .aout3(aout27_8), .aout4(aout28_8),
                    .wout1(wout28_5), .wout2(wout28_6), .wout3(wout28_7), .wout4(wout28_8),
                    .sout11(sout25_5), .sout12(sout25_6), .sout13(sout25_7), .sout14(sout25_8),
                    .sout21(sout26_5), .sout22(sout26_6), .sout23(sout26_7), .sout24(sout26_8),
                    .sout31(sout27_5), .sout32(sout27_6), .sout33(sout27_7), .sout34(sout27_8),
                    .sout41(sout28_5), .sout42(sout28_6), .sout43(sout28_7), .sout44(sout28_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_73 (.clk(clk), .rst(rst),
                    .ain1(aout25_8), .ain2(aout26_8), .ain3(aout27_8), .ain4(aout28_8),
                    .win1(wout24_9), .win2(wout24_10), .win3(wout24_11), .win4(wout24_12),
                    .aout1(aout25_12), .aout2(aout26_12), .aout3(aout27_12), .aout4(aout28_12),
                    .wout1(wout28_9), .wout2(wout28_10), .wout3(wout28_11), .wout4(wout28_12),
                    .sout11(sout25_9), .sout12(sout25_10), .sout13(sout25_11), .sout14(sout25_12),
                    .sout21(sout26_9), .sout22(sout26_10), .sout23(sout26_11), .sout24(sout26_12),
                    .sout31(sout27_9), .sout32(sout27_10), .sout33(sout27_11), .sout34(sout27_12),
                    .sout41(sout28_9), .sout42(sout28_10), .sout43(sout28_11), .sout44(sout28_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_74 (.clk(clk), .rst(rst),
                    .ain1(aout25_12), .ain2(aout26_12), .ain3(aout27_12), .ain4(aout28_12),
                    .win1(wout24_13), .win2(wout24_14), .win3(wout24_15), .win4(wout24_16),
                    .aout1(aout25_16), .aout2(aout26_16), .aout3(aout27_16), .aout4(aout28_16),
                    .wout1(wout28_13), .wout2(wout28_14), .wout3(wout28_15), .wout4(wout28_16),
                    .sout11(sout25_13), .sout12(sout25_14), .sout13(sout25_15), .sout14(sout25_16),
                    .sout21(sout26_13), .sout22(sout26_14), .sout23(sout26_15), .sout24(sout26_16),
                    .sout31(sout27_13), .sout32(sout27_14), .sout33(sout27_15), .sout34(sout27_16),
                    .sout41(sout28_13), .sout42(sout28_14), .sout43(sout28_15), .sout44(sout28_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_75 (.clk(clk), .rst(rst),
                    .ain1(aout25_16), .ain2(aout26_16), .ain3(aout27_16), .ain4(aout28_16),
                    .win1(wout24_17), .win2(wout24_18), .win3(wout24_19), .win4(wout24_20),
                    .aout1(aout25_20), .aout2(aout26_20), .aout3(aout27_20), .aout4(aout28_20),
                    .wout1(wout28_17), .wout2(wout28_18), .wout3(wout28_19), .wout4(wout28_20),
                    .sout11(sout25_17), .sout12(sout25_18), .sout13(sout25_19), .sout14(sout25_20),
                    .sout21(sout26_17), .sout22(sout26_18), .sout23(sout26_19), .sout24(sout26_20),
                    .sout31(sout27_17), .sout32(sout27_18), .sout33(sout27_19), .sout34(sout27_20),
                    .sout41(sout28_17), .sout42(sout28_18), .sout43(sout28_19), .sout44(sout28_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_76 (.clk(clk), .rst(rst),
                    .ain1(aout25_20), .ain2(aout26_20), .ain3(aout27_20), .ain4(aout28_20),
                    .win1(wout24_21), .win2(wout24_22), .win3(wout24_23), .win4(wout24_24),
                    .aout1(aout25_24), .aout2(aout26_24), .aout3(aout27_24), .aout4(aout28_24),
                    .wout1(wout28_21), .wout2(wout28_22), .wout3(wout28_23), .wout4(wout28_24),
                    .sout11(sout25_21), .sout12(sout25_22), .sout13(sout25_23), .sout14(sout25_24),
                    .sout21(sout26_21), .sout22(sout26_22), .sout23(sout26_23), .sout24(sout26_24),
                    .sout31(sout27_21), .sout32(sout27_22), .sout33(sout27_23), .sout34(sout27_24),
                    .sout41(sout28_21), .sout42(sout28_22), .sout43(sout28_23), .sout44(sout28_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_77 (.clk(clk), .rst(rst),
                    .ain1(aout25_24), .ain2(aout26_24), .ain3(aout27_24), .ain4(aout28_24),
                    .win1(wout24_25), .win2(wout24_26), .win3(wout24_27), .win4(wout24_28),
                    .aout1(aout25_28), .aout2(aout26_28), .aout3(aout27_28), .aout4(aout28_28),
                    .wout1(wout28_25), .wout2(wout28_26), .wout3(wout28_27), .wout4(wout28_28),
                    .sout11(sout25_25), .sout12(sout25_26), .sout13(sout25_27), .sout14(sout25_28),
                    .sout21(sout26_25), .sout22(sout26_26), .sout23(sout26_27), .sout24(sout26_28),
                    .sout31(sout27_25), .sout32(sout27_26), .sout33(sout27_27), .sout34(sout27_28),
                    .sout41(sout28_25), .sout42(sout28_26), .sout43(sout28_27), .sout44(sout28_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_78 (.clk(clk), .rst(rst),
                    .ain1(aout25_28), .ain2(aout26_28), .ain3(aout27_28), .ain4(aout28_28),
                    .win1(wout24_29), .win2(wout24_30), .win3(wout24_31), .win4(wout24_32),
                    .aout1(aout25_32), .aout2(aout26_32), .aout3(aout27_32), .aout4(aout28_32),
                    .wout1(wout28_29), .wout2(wout28_30), .wout3(wout28_31), .wout4(wout28_32),
                    .sout11(sout25_29), .sout12(sout25_30), .sout13(sout25_31), .sout14(sout25_32),
                    .sout21(sout26_29), .sout22(sout26_30), .sout23(sout26_31), .sout24(sout26_32),
                    .sout31(sout27_29), .sout32(sout27_30), .sout33(sout27_31), .sout34(sout27_32),
                    .sout41(sout28_29), .sout42(sout28_30), .sout43(sout28_31), .sout44(sout28_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_79 (.clk(clk), .rst(rst),
                    .ain1(aout25_32), .ain2(aout26_32), .ain3(aout27_32), .ain4(aout28_32),
                    .win1(wout24_33), .win2(wout24_34), .win3(wout24_35), .win4(wout24_36),
                    .aout1(aout25_36), .aout2(aout26_36), .aout3(aout27_36), .aout4(aout28_36),
                    .wout1(wout28_33), .wout2(wout28_34), .wout3(wout28_35), .wout4(wout28_36),
                    .sout11(sout25_33), .sout12(sout25_34), .sout13(sout25_35), .sout14(sout25_36),
                    .sout21(sout26_33), .sout22(sout26_34), .sout23(sout26_35), .sout24(sout26_36),
                    .sout31(sout27_33), .sout32(sout27_34), .sout33(sout27_35), .sout34(sout27_36),
                    .sout41(sout28_33), .sout42(sout28_34), .sout43(sout28_35), .sout44(sout28_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_7_10 (.clk(clk), .rst(rst),
                    .ain1(aout25_36), .ain2(aout26_36), .ain3(aout27_36), .ain4(aout28_36),
                    .win1(wout24_37), .win2(wout24_38), .win3(wout24_39), .win4(wout24_40),
                    .aout1(aout25_40), .aout2(aout26_40), .aout3(aout27_40), .aout4(aout28_40),
                    .wout1(wout28_37), .wout2(wout28_38), .wout3(wout28_39), .wout4(wout28_40),
                    .sout11(sout25_37), .sout12(sout25_38), .sout13(sout25_39), .sout14(sout25_40),
                    .sout21(sout26_37), .sout22(sout26_38), .sout23(sout26_39), .sout24(sout26_40),
                    .sout31(sout27_37), .sout32(sout27_38), .sout33(sout27_39), .sout34(sout27_40),
                    .sout41(sout28_37), .sout42(sout28_38), .sout43(sout28_39), .sout44(sout28_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_7_11 (.clk(clk), .rst(rst),
                    .ain1(aout25_40), .ain2(aout26_40), .ain3(aout27_40), .ain4(aout28_40),
                    .win1(wout24_41), .win2(wout24_42), .win3(wout24_43), .win4(wout24_44),
                    .aout1(aout25_44), .aout2(aout26_44), .aout3(aout27_44), .aout4(aout28_44),
                    .wout1(wout28_41), .wout2(wout28_42), .wout3(wout28_43), .wout4(wout28_44),
                    .sout11(sout25_41), .sout12(sout25_42), .sout13(sout25_43), .sout14(sout25_44),
                    .sout21(sout26_41), .sout22(sout26_42), .sout23(sout26_43), .sout24(sout26_44),
                    .sout31(sout27_41), .sout32(sout27_42), .sout33(sout27_43), .sout34(sout27_44),
                    .sout41(sout28_41), .sout42(sout28_42), .sout43(sout28_43), .sout44(sout28_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_7_12 (.clk(clk), .rst(rst),
                    .ain1(aout25_44), .ain2(aout26_44), .ain3(aout27_44), .ain4(aout28_44),
                    .win1(wout24_45), .win2(wout24_46), .win3(wout24_47), .win4(wout24_48),
                    .aout1(aout25_48), .aout2(aout26_48), .aout3(aout27_48), .aout4(aout28_48),
                    .wout1(wout28_45), .wout2(wout28_46), .wout3(wout28_47), .wout4(wout28_48),
                    .sout11(sout25_45), .sout12(sout25_46), .sout13(sout25_47), .sout14(sout25_48),
                    .sout21(sout26_45), .sout22(sout26_46), .sout23(sout26_47), .sout24(sout26_48),
                    .sout31(sout27_45), .sout32(sout27_46), .sout33(sout27_47), .sout34(sout27_48),
                    .sout41(sout28_45), .sout42(sout28_46), .sout43(sout28_47), .sout44(sout28_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_7_13 (.clk(clk), .rst(rst),
                    .ain1(aout25_48), .ain2(aout26_48), .ain3(aout27_48), .ain4(aout28_48),
                    .win1(wout24_49), .win2(wout24_50), .win3(wout24_51), .win4(wout24_52),
                    .aout1(aout25_52), .aout2(aout26_52), .aout3(aout27_52), .aout4(aout28_52),
                    .wout1(wout28_49), .wout2(wout28_50), .wout3(wout28_51), .wout4(wout28_52),
                    .sout11(sout25_49), .sout12(sout25_50), .sout13(sout25_51), .sout14(sout25_52),
                    .sout21(sout26_49), .sout22(sout26_50), .sout23(sout26_51), .sout24(sout26_52),
                    .sout31(sout27_49), .sout32(sout27_50), .sout33(sout27_51), .sout34(sout27_52),
                    .sout41(sout28_49), .sout42(sout28_50), .sout43(sout28_51), .sout44(sout28_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_7_14 (.clk(clk), .rst(rst),
                    .ain1(aout25_52), .ain2(aout26_52), .ain3(aout27_52), .ain4(aout28_52),
                    .win1(wout24_53), .win2(wout24_54), .win3(wout24_55), .win4(wout24_56),
                    .aout1(aout25_56), .aout2(aout26_56), .aout3(aout27_56), .aout4(aout28_56),
                    .wout1(wout28_53), .wout2(wout28_54), .wout3(wout28_55), .wout4(wout28_56),
                    .sout11(sout25_53), .sout12(sout25_54), .sout13(sout25_55), .sout14(sout25_56),
                    .sout21(sout26_53), .sout22(sout26_54), .sout23(sout26_55), .sout24(sout26_56),
                    .sout31(sout27_53), .sout32(sout27_54), .sout33(sout27_55), .sout34(sout27_56),
                    .sout41(sout28_53), .sout42(sout28_54), .sout43(sout28_55), .sout44(sout28_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_7_15 (.clk(clk), .rst(rst),
                    .ain1(aout25_56), .ain2(aout26_56), .ain3(aout27_56), .ain4(aout28_56),
                    .win1(wout24_57), .win2(wout24_58), .win3(wout24_59), .win4(wout24_60),
                    .aout1(aout25_60), .aout2(aout26_60), .aout3(aout27_60), .aout4(aout28_60),
                    .wout1(wout28_57), .wout2(wout28_58), .wout3(wout28_59), .wout4(wout28_60),
                    .sout11(sout25_57), .sout12(sout25_58), .sout13(sout25_59), .sout14(sout25_60),
                    .sout21(sout26_57), .sout22(sout26_58), .sout23(sout26_59), .sout24(sout26_60),
                    .sout31(sout27_57), .sout32(sout27_58), .sout33(sout27_59), .sout34(sout27_60),
                    .sout41(sout28_57), .sout42(sout28_58), .sout43(sout28_59), .sout44(sout28_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_7_16 (.clk(clk), .rst(rst),
                    .ain1(aout25_60), .ain2(aout26_60), .ain3(aout27_60), .ain4(aout28_60),
                    .win1(wout24_61), .win2(wout24_62), .win3(wout24_63), .win4(wout24_64),
                    .aout1(aout25_64), .aout2(aout26_64), .aout3(aout27_64), .aout4(aout28_64),
                    .wout1(wout28_61), .wout2(wout28_62), .wout3(wout28_63), .wout4(wout28_64),
                    .sout11(sout25_61), .sout12(sout25_62), .sout13(sout25_63), .sout14(sout25_64),
                    .sout21(sout26_61), .sout22(sout26_62), .sout23(sout26_63), .sout24(sout26_64),
                    .sout31(sout27_61), .sout32(sout27_62), .sout33(sout27_63), .sout34(sout27_64),
                    .sout41(sout28_61), .sout42(sout28_62), .sout43(sout28_63), .sout44(sout28_64)
                    ); //4x4 MAC array
    
    //row8    
    mac_array_4x4 mac_array_4x4_81 (.clk(clk), .rst(rst),
                    .ain1(ain29), .ain2(ain30), .ain3(ain31), .ain4(ain32),
                    .win1(wout28_1), .win2(wout28_2), .win3(wout28_3), .win4(wout28_4),
                    .aout1(aout29_4), .aout2(aout30_4), .aout3(aout31_4), .aout4(aout32_4),
                    .wout1(wout32_1), .wout2(wout32_2), .wout3(wout32_3), .wout4(wout32_4),
                    .sout11(sout29_1), .sout12(sout29_2), .sout13(sout29_3), .sout14(sout29_4),
                    .sout21(sout30_1), .sout22(sout30_2), .sout23(sout30_3), .sout24(sout30_4),
                    .sout31(sout31_1), .sout32(sout31_2), .sout33(sout31_3), .sout34(sout31_4),
                    .sout41(sout32_1), .sout42(sout32_2), .sout43(sout32_3), .sout44(sout32_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_82 (.clk(clk), .rst(rst),
                    .ain1(aout29_4), .ain2(aout30_4), .ain3(aout31_4), .ain4(aout32_4),
                    .win1(wout28_5), .win2(wout28_6), .win3(wout28_7), .win4(wout28_8),
                    .aout1(aout29_8), .aout2(aout30_8), .aout3(aout31_8), .aout4(aout32_8),
                    .wout1(wout32_5), .wout2(wout32_6), .wout3(wout32_7), .wout4(wout32_8),
                    .sout11(sout29_5), .sout12(sout29_6), .sout13(sout29_7), .sout14(sout29_8),
                    .sout21(sout30_5), .sout22(sout30_6), .sout23(sout30_7), .sout24(sout30_8),
                    .sout31(sout31_5), .sout32(sout31_6), .sout33(sout31_7), .sout34(sout31_8),
                    .sout41(sout32_5), .sout42(sout32_6), .sout43(sout32_7), .sout44(sout32_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_83 (.clk(clk), .rst(rst),
                    .ain1(aout29_8), .ain2(aout30_8), .ain3(aout31_8), .ain4(aout32_8),
                    .win1(wout28_9), .win2(wout28_10), .win3(wout28_11), .win4(wout28_12),
                    .aout1(aout29_12), .aout2(aout30_12), .aout3(aout31_12), .aout4(aout32_12),
                    .wout1(wout32_9), .wout2(wout32_10), .wout3(wout32_11), .wout4(wout32_12),
                    .sout11(sout29_9), .sout12(sout29_10), .sout13(sout29_11), .sout14(sout29_12),
                    .sout21(sout30_9), .sout22(sout30_10), .sout23(sout30_11), .sout24(sout30_12),
                    .sout31(sout31_9), .sout32(sout31_10), .sout33(sout31_11), .sout34(sout31_12),
                    .sout41(sout32_9), .sout42(sout32_10), .sout43(sout32_11), .sout44(sout32_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_84 (.clk(clk), .rst(rst),
                    .ain1(aout29_12), .ain2(aout30_12), .ain3(aout31_12), .ain4(aout32_12),
                    .win1(wout28_13), .win2(wout28_14), .win3(wout28_15), .win4(wout28_16),
                    .aout1(aout29_16), .aout2(aout30_16), .aout3(aout31_16), .aout4(aout32_16),
                    .wout1(wout32_13), .wout2(wout32_14), .wout3(wout32_15), .wout4(wout32_16),
                    .sout11(sout29_13), .sout12(sout29_14), .sout13(sout29_15), .sout14(sout29_16),
                    .sout21(sout30_13), .sout22(sout30_14), .sout23(sout30_15), .sout24(sout30_16),
                    .sout31(sout31_13), .sout32(sout31_14), .sout33(sout31_15), .sout34(sout31_16),
                    .sout41(sout32_13), .sout42(sout32_14), .sout43(sout32_15), .sout44(sout32_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_85 (.clk(clk), .rst(rst),
                    .ain1(aout29_16), .ain2(aout30_16), .ain3(aout31_16), .ain4(aout32_16),
                    .win1(wout28_17), .win2(wout28_18), .win3(wout28_19), .win4(wout28_20),
                    .aout1(aout29_20), .aout2(aout30_20), .aout3(aout31_20), .aout4(aout32_20),
                    .wout1(wout32_17), .wout2(wout32_18), .wout3(wout32_19), .wout4(wout32_20),
                    .sout11(sout29_17), .sout12(sout29_18), .sout13(sout29_19), .sout14(sout29_20),
                    .sout21(sout30_17), .sout22(sout30_18), .sout23(sout30_19), .sout24(sout30_20),
                    .sout31(sout31_17), .sout32(sout31_18), .sout33(sout31_19), .sout34(sout31_20),
                    .sout41(sout32_17), .sout42(sout32_18), .sout43(sout32_19), .sout44(sout32_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_86 (.clk(clk), .rst(rst),
                    .ain1(aout29_20), .ain2(aout30_20), .ain3(aout31_20), .ain4(aout32_20),
                    .win1(wout28_21), .win2(wout28_22), .win3(wout28_23), .win4(wout28_24),
                    .aout1(aout29_24), .aout2(aout30_24), .aout3(aout31_24), .aout4(aout32_24),
                    .wout1(wout32_21), .wout2(wout32_22), .wout3(wout32_23), .wout4(wout32_24),
                    .sout11(sout29_21), .sout12(sout29_22), .sout13(sout29_23), .sout14(sout29_24),
                    .sout21(sout30_21), .sout22(sout30_22), .sout23(sout30_23), .sout24(sout30_24),
                    .sout31(sout31_21), .sout32(sout31_22), .sout33(sout31_23), .sout34(sout31_24),
                    .sout41(sout32_21), .sout42(sout32_22), .sout43(sout32_23), .sout44(sout32_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_87 (.clk(clk), .rst(rst),
                    .ain1(aout29_24), .ain2(aout30_24), .ain3(aout31_24), .ain4(aout32_24),
                    .win1(wout28_25), .win2(wout28_26), .win3(wout28_27), .win4(wout28_28),
                    .aout1(aout29_28), .aout2(aout30_28), .aout3(aout31_28), .aout4(aout32_28),
                    .wout1(wout32_25), .wout2(wout32_26), .wout3(wout32_27), .wout4(wout32_28),
                    .sout11(sout29_25), .sout12(sout29_26), .sout13(sout29_27), .sout14(sout29_28),
                    .sout21(sout30_25), .sout22(sout30_26), .sout23(sout30_27), .sout24(sout30_28),
                    .sout31(sout31_25), .sout32(sout31_26), .sout33(sout31_27), .sout34(sout31_28),
                    .sout41(sout32_25), .sout42(sout32_26), .sout43(sout32_27), .sout44(sout32_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_88 (.clk(clk), .rst(rst),
                    .ain1(aout29_28), .ain2(aout30_28), .ain3(aout31_28), .ain4(aout32_28),
                    .win1(wout28_29), .win2(wout28_30), .win3(wout28_31), .win4(wout28_32),
                    .aout1(aout29_32), .aout2(aout30_32), .aout3(aout31_32), .aout4(aout32_32),
                    .wout1(wout32_29), .wout2(wout32_30), .wout3(wout32_31), .wout4(wout32_32),
                    .sout11(sout29_29), .sout12(sout29_30), .sout13(sout29_31), .sout14(sout29_32),
                    .sout21(sout30_29), .sout22(sout30_30), .sout23(sout30_31), .sout24(sout30_32),
                    .sout31(sout31_29), .sout32(sout31_30), .sout33(sout31_31), .sout34(sout31_32),
                    .sout41(sout32_29), .sout42(sout32_30), .sout43(sout32_31), .sout44(sout32_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_89 (.clk(clk), .rst(rst),
                    .ain1(aout29_32), .ain2(aout30_32), .ain3(aout31_32), .ain4(aout32_32),
                    .win1(wout28_33), .win2(wout28_34), .win3(wout28_35), .win4(wout28_36),
                    .aout1(aout29_36), .aout2(aout30_36), .aout3(aout31_36), .aout4(aout32_36),
                    .wout1(wout32_33), .wout2(wout32_34), .wout3(wout32_35), .wout4(wout32_36),
                    .sout11(sout29_33), .sout12(sout29_34), .sout13(sout29_35), .sout14(sout29_36),
                    .sout21(sout30_33), .sout22(sout30_34), .sout23(sout30_35), .sout24(sout30_36),
                    .sout31(sout31_33), .sout32(sout31_34), .sout33(sout31_35), .sout34(sout31_36),
                    .sout41(sout32_33), .sout42(sout32_34), .sout43(sout32_35), .sout44(sout32_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_8_10 (.clk(clk), .rst(rst),
                    .ain1(aout29_36), .ain2(aout30_36), .ain3(aout31_36), .ain4(aout32_36),
                    .win1(wout28_37), .win2(wout28_38), .win3(wout28_39), .win4(wout28_40),
                    .aout1(aout29_40), .aout2(aout30_40), .aout3(aout31_40), .aout4(aout32_40),
                    .wout1(wout32_37), .wout2(wout32_38), .wout3(wout32_39), .wout4(wout32_40),
                    .sout11(sout29_37), .sout12(sout29_38), .sout13(sout29_39), .sout14(sout29_40),
                    .sout21(sout30_37), .sout22(sout30_38), .sout23(sout30_39), .sout24(sout30_40),
                    .sout31(sout31_37), .sout32(sout31_38), .sout33(sout31_39), .sout34(sout31_40),
                    .sout41(sout32_37), .sout42(sout32_38), .sout43(sout32_39), .sout44(sout32_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_8_11 (.clk(clk), .rst(rst),
                    .ain1(aout29_40), .ain2(aout30_40), .ain3(aout31_40), .ain4(aout32_40),
                    .win1(wout28_41), .win2(wout28_42), .win3(wout28_43), .win4(wout28_44),
                    .aout1(aout29_44), .aout2(aout30_44), .aout3(aout31_44), .aout4(aout32_44),
                    .wout1(wout32_41), .wout2(wout32_42), .wout3(wout32_43), .wout4(wout32_44),
                    .sout11(sout29_41), .sout12(sout29_42), .sout13(sout29_43), .sout14(sout29_44),
                    .sout21(sout30_41), .sout22(sout30_42), .sout23(sout30_43), .sout24(sout30_44),
                    .sout31(sout31_41), .sout32(sout31_42), .sout33(sout31_43), .sout34(sout31_44),
                    .sout41(sout32_41), .sout42(sout32_42), .sout43(sout32_43), .sout44(sout32_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_8_12 (.clk(clk), .rst(rst),
                    .ain1(aout29_44), .ain2(aout30_44), .ain3(aout31_44), .ain4(aout32_44),
                    .win1(wout28_45), .win2(wout28_46), .win3(wout28_47), .win4(wout28_48),
                    .aout1(aout29_48), .aout2(aout30_48), .aout3(aout31_48), .aout4(aout32_48),
                    .wout1(wout32_45), .wout2(wout32_46), .wout3(wout32_47), .wout4(wout32_48),
                    .sout11(sout29_45), .sout12(sout29_46), .sout13(sout29_47), .sout14(sout29_48),
                    .sout21(sout30_45), .sout22(sout30_46), .sout23(sout30_47), .sout24(sout30_48),
                    .sout31(sout31_45), .sout32(sout31_46), .sout33(sout31_47), .sout34(sout31_48),
                    .sout41(sout32_45), .sout42(sout32_46), .sout43(sout32_47), .sout44(sout32_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_8_13 (.clk(clk), .rst(rst),
                    .ain1(aout29_48), .ain2(aout30_48), .ain3(aout31_48), .ain4(aout32_48),
                    .win1(wout28_49), .win2(wout28_50), .win3(wout28_51), .win4(wout28_52),
                    .aout1(aout29_52), .aout2(aout30_52), .aout3(aout31_52), .aout4(aout32_52),
                    .wout1(wout32_49), .wout2(wout32_50), .wout3(wout32_51), .wout4(wout32_52),
                    .sout11(sout29_49), .sout12(sout29_50), .sout13(sout29_51), .sout14(sout29_52),
                    .sout21(sout30_49), .sout22(sout30_50), .sout23(sout30_51), .sout24(sout30_52),
                    .sout31(sout31_49), .sout32(sout31_50), .sout33(sout31_51), .sout34(sout31_52),
                    .sout41(sout32_49), .sout42(sout32_50), .sout43(sout32_51), .sout44(sout32_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_8_14 (.clk(clk), .rst(rst),
                    .ain1(aout29_52), .ain2(aout30_52), .ain3(aout31_52), .ain4(aout32_52),
                    .win1(wout28_53), .win2(wout28_54), .win3(wout28_55), .win4(wout28_56),
                    .aout1(aout29_56), .aout2(aout30_56), .aout3(aout31_56), .aout4(aout32_56),
                    .wout1(wout32_53), .wout2(wout32_54), .wout3(wout32_55), .wout4(wout32_56),
                    .sout11(sout29_53), .sout12(sout29_54), .sout13(sout29_55), .sout14(sout29_56),
                    .sout21(sout30_53), .sout22(sout30_54), .sout23(sout30_55), .sout24(sout30_56),
                    .sout31(sout31_53), .sout32(sout31_54), .sout33(sout31_55), .sout34(sout31_56),
                    .sout41(sout32_53), .sout42(sout32_54), .sout43(sout32_55), .sout44(sout32_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_8_15 (.clk(clk), .rst(rst),
                    .ain1(aout29_56), .ain2(aout30_56), .ain3(aout31_56), .ain4(aout32_56),
                    .win1(wout28_57), .win2(wout28_58), .win3(wout28_59), .win4(wout28_60),
                    .aout1(aout29_60), .aout2(aout30_60), .aout3(aout31_60), .aout4(aout32_60),
                    .wout1(wout32_57), .wout2(wout32_58), .wout3(wout32_59), .wout4(wout32_60),
                    .sout11(sout29_57), .sout12(sout29_58), .sout13(sout29_59), .sout14(sout29_60),
                    .sout21(sout30_57), .sout22(sout30_58), .sout23(sout30_59), .sout24(sout30_60),
                    .sout31(sout31_57), .sout32(sout31_58), .sout33(sout31_59), .sout34(sout31_60),
                    .sout41(sout32_57), .sout42(sout32_58), .sout43(sout32_59), .sout44(sout32_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_8_16 (.clk(clk), .rst(rst),
                    .ain1(aout29_60), .ain2(aout30_60), .ain3(aout31_60), .ain4(aout32_60),
                    .win1(wout28_61), .win2(wout28_62), .win3(wout28_63), .win4(wout28_64),
                    .aout1(aout29_64), .aout2(aout30_64), .aout3(aout31_64), .aout4(aout32_64),
                    .wout1(wout32_61), .wout2(wout32_62), .wout3(wout32_63), .wout4(wout32_64),
                    .sout11(sout29_61), .sout12(sout29_62), .sout13(sout29_63), .sout14(sout29_64),
                    .sout21(sout30_61), .sout22(sout30_62), .sout23(sout30_63), .sout24(sout30_64),
                    .sout31(sout31_61), .sout32(sout31_62), .sout33(sout31_63), .sout34(sout31_64),
                    .sout41(sout32_61), .sout42(sout32_62), .sout43(sout32_63), .sout44(sout32_64)
                    ); //4x4 MAC array
                    
  
    //row9   
    mac_array_4x4 mac_array_4x4_91 (.clk(clk), .rst(rst),
                    .ain1(ain33), .ain2(ain34), .ain3(ain35), .ain4(ain36),
                    .win1(wout32_1), .win2(wout32_2), .win3(wout32_3), .win4(wout32_4),
                    .aout1(aout33_4), .aout2(aout34_4), .aout3(aout35_4), .aout4(aout36_4),
                    .wout1(wout36_1), .wout2(wout36_2), .wout3(wout36_3), .wout4(wout36_4),
                    .sout11(sout33_1), .sout12(sout33_2), .sout13(sout33_3), .sout14(sout33_4),
                    .sout21(sout34_1), .sout22(sout34_2), .sout23(sout34_3), .sout24(sout34_4),
                    .sout31(sout35_1), .sout32(sout35_2), .sout33(sout35_3), .sout34(sout35_4),
                    .sout41(sout36_1), .sout42(sout36_2), .sout43(sout36_3), .sout44(sout36_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_92 (.clk(clk), .rst(rst),
                    .ain1(aout33_4), .ain2(aout34_4), .ain3(aout35_4), .ain4(aout36_4),
                    .win1(wout32_5), .win2(wout32_6), .win3(wout32_7), .win4(wout32_8),
                    .aout1(aout33_8), .aout2(aout34_8), .aout3(aout35_8), .aout4(aout36_8),
                    .wout1(wout36_5), .wout2(wout36_6), .wout3(wout36_7), .wout4(wout36_8),
                    .sout11(sout33_5), .sout12(sout33_6), .sout13(sout33_7), .sout14(sout33_8),
                    .sout21(sout34_5), .sout22(sout34_6), .sout23(sout34_7), .sout24(sout34_8),
                    .sout31(sout35_5), .sout32(sout35_6), .sout33(sout35_7), .sout34(sout35_8),
                    .sout41(sout36_5), .sout42(sout36_6), .sout43(sout36_7), .sout44(sout36_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_93 (.clk(clk), .rst(rst),
                    .ain1(aout33_8), .ain2(aout34_8), .ain3(aout35_8), .ain4(aout36_8),
                    .win1(wout32_9), .win2(wout32_10), .win3(wout32_11), .win4(wout32_12),
                    .aout1(aout33_12), .aout2(aout34_12), .aout3(aout35_12), .aout4(aout36_12),
                    .wout1(wout36_9), .wout2(wout36_10), .wout3(wout36_11), .wout4(wout36_12),
                    .sout11(sout33_9), .sout12(sout33_10), .sout13(sout33_11), .sout14(sout33_12),
                    .sout21(sout34_9), .sout22(sout34_10), .sout23(sout34_11), .sout24(sout34_12),
                    .sout31(sout35_9), .sout32(sout35_10), .sout33(sout35_11), .sout34(sout35_12),
                    .sout41(sout36_9), .sout42(sout36_10), .sout43(sout36_11), .sout44(sout36_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_94 (.clk(clk), .rst(rst),
                    .ain1(aout33_12), .ain2(aout34_12), .ain3(aout35_12), .ain4(aout36_12),
                    .win1(wout32_13), .win2(wout32_14), .win3(wout32_15), .win4(wout32_16),
                    .aout1(aout33_16), .aout2(aout34_16), .aout3(aout35_16), .aout4(aout36_16),
                    .wout1(wout36_13), .wout2(wout36_14), .wout3(wout36_15), .wout4(wout36_16),
                    .sout11(sout33_13), .sout12(sout33_14), .sout13(sout33_15), .sout14(sout33_16),
                    .sout21(sout34_13), .sout22(sout34_14), .sout23(sout34_15), .sout24(sout34_16),
                    .sout31(sout35_13), .sout32(sout35_14), .sout33(sout35_15), .sout34(sout35_16),
                    .sout41(sout36_13), .sout42(sout36_14), .sout43(sout36_15), .sout44(sout36_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_95 (.clk(clk), .rst(rst),
                    .ain1(aout33_16), .ain2(aout34_16), .ain3(aout35_16), .ain4(aout36_16),
                    .win1(wout32_17), .win2(wout32_18), .win3(wout32_19), .win4(wout32_20),
                    .aout1(aout33_20), .aout2(aout34_20), .aout3(aout35_20), .aout4(aout36_20),
                    .wout1(wout36_17), .wout2(wout36_18), .wout3(wout36_19), .wout4(wout36_20),
                    .sout11(sout33_17), .sout12(sout33_18), .sout13(sout33_19), .sout14(sout33_20),
                    .sout21(sout34_17), .sout22(sout34_18), .sout23(sout34_19), .sout24(sout34_20),
                    .sout31(sout35_17), .sout32(sout35_18), .sout33(sout35_19), .sout34(sout35_20),
                    .sout41(sout36_17), .sout42(sout36_18), .sout43(sout36_19), .sout44(sout36_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_96 (.clk(clk), .rst(rst),
                    .ain1(aout33_20), .ain2(aout34_20), .ain3(aout35_20), .ain4(aout36_20),
                    .win1(wout32_21), .win2(wout32_22), .win3(wout32_23), .win4(wout32_24),
                    .aout1(aout33_24), .aout2(aout34_24), .aout3(aout35_24), .aout4(aout36_24),
                    .wout1(wout36_21), .wout2(wout36_22), .wout3(wout36_23), .wout4(wout36_24),
                    .sout11(sout33_21), .sout12(sout33_22), .sout13(sout33_23), .sout14(sout33_24),
                    .sout21(sout34_21), .sout22(sout34_22), .sout23(sout34_23), .sout24(sout34_24),
                    .sout31(sout35_21), .sout32(sout35_22), .sout33(sout35_23), .sout34(sout35_24),
                    .sout41(sout36_21), .sout42(sout36_22), .sout43(sout36_23), .sout44(sout36_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_97 (.clk(clk), .rst(rst),
                    .ain1(aout33_24), .ain2(aout34_24), .ain3(aout35_24), .ain4(aout36_24),
                    .win1(wout32_25), .win2(wout32_26), .win3(wout32_27), .win4(wout32_28),
                    .aout1(aout33_28), .aout2(aout34_28), .aout3(aout35_28), .aout4(aout36_28),
                    .wout1(wout36_25), .wout2(wout36_26), .wout3(wout36_27), .wout4(wout36_28),
                    .sout11(sout33_25), .sout12(sout33_26), .sout13(sout33_27), .sout14(sout33_28),
                    .sout21(sout34_25), .sout22(sout34_26), .sout23(sout34_27), .sout24(sout34_28),
                    .sout31(sout35_25), .sout32(sout35_26), .sout33(sout35_27), .sout34(sout35_28),
                    .sout41(sout36_25), .sout42(sout36_26), .sout43(sout36_27), .sout44(sout36_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_98 (.clk(clk), .rst(rst),
                    .ain1(aout33_28), .ain2(aout34_28), .ain3(aout35_28), .ain4(aout36_28),
                    .win1(wout32_29), .win2(wout32_30), .win3(wout32_31), .win4(wout32_32),
                    .aout1(aout33_32), .aout2(aout34_32), .aout3(aout35_32), .aout4(aout36_32),
                    .wout1(wout36_29), .wout2(wout36_30), .wout3(wout36_31), .wout4(wout36_32),
                    .sout11(sout33_29), .sout12(sout33_30), .sout13(sout33_31), .sout14(sout33_32),
                    .sout21(sout34_29), .sout22(sout34_30), .sout23(sout34_31), .sout24(sout34_32),
                    .sout31(sout35_29), .sout32(sout35_30), .sout33(sout35_31), .sout34(sout35_32),
                    .sout41(sout36_29), .sout42(sout36_30), .sout43(sout36_31), .sout44(sout36_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_99 (.clk(clk), .rst(rst),
                    .ain1(aout33_32), .ain2(aout34_32), .ain3(aout35_32), .ain4(aout36_32),
                    .win1(wout32_33), .win2(wout32_34), .win3(wout32_35), .win4(wout32_36),
                    .aout1(aout33_36), .aout2(aout34_36), .aout3(aout35_36), .aout4(aout36_36),
                    .wout1(wout36_33), .wout2(wout36_34), .wout3(wout36_35), .wout4(wout36_36),
                    .sout11(sout33_33), .sout12(sout33_34), .sout13(sout33_35), .sout14(sout33_36),
                    .sout21(sout34_33), .sout22(sout34_34), .sout23(sout34_35), .sout24(sout34_36),
                    .sout31(sout35_33), .sout32(sout35_34), .sout33(sout35_35), .sout34(sout35_36),
                    .sout41(sout36_33), .sout42(sout36_34), .sout43(sout36_35), .sout44(sout36_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_9_10 (.clk(clk), .rst(rst),
                    .ain1(aout33_36), .ain2(aout34_36), .ain3(aout35_36), .ain4(aout36_36),
                    .win1(wout32_37), .win2(wout32_38), .win3(wout32_39), .win4(wout32_40),
                    .aout1(aout33_40), .aout2(aout34_40), .aout3(aout35_40), .aout4(aout36_40),
                    .wout1(wout36_37), .wout2(wout36_38), .wout3(wout36_39), .wout4(wout36_40),
                    .sout11(sout33_37), .sout12(sout33_38), .sout13(sout33_39), .sout14(sout33_40),
                    .sout21(sout34_37), .sout22(sout34_38), .sout23(sout34_39), .sout24(sout34_40),
                    .sout31(sout35_37), .sout32(sout35_38), .sout33(sout35_39), .sout34(sout35_40),
                    .sout41(sout36_37), .sout42(sout36_38), .sout43(sout36_39), .sout44(sout36_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_9_11 (.clk(clk), .rst(rst),
                    .ain1(aout33_40), .ain2(aout34_40), .ain3(aout35_40), .ain4(aout36_40),
                    .win1(wout32_41), .win2(wout32_42), .win3(wout32_43), .win4(wout32_44),
                    .aout1(aout33_44), .aout2(aout34_44), .aout3(aout35_44), .aout4(aout36_44),
                    .wout1(wout36_41), .wout2(wout36_42), .wout3(wout36_43), .wout4(wout36_44),
                    .sout11(sout33_41), .sout12(sout33_42), .sout13(sout33_43), .sout14(sout33_44),
                    .sout21(sout34_41), .sout22(sout34_42), .sout23(sout34_43), .sout24(sout34_44),
                    .sout31(sout35_41), .sout32(sout35_42), .sout33(sout35_43), .sout34(sout35_44),
                    .sout41(sout36_41), .sout42(sout36_42), .sout43(sout36_43), .sout44(sout36_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_9_12 (.clk(clk), .rst(rst),
                    .ain1(aout33_44), .ain2(aout34_44), .ain3(aout35_44), .ain4(aout36_44),
                    .win1(wout32_45), .win2(wout32_46), .win3(wout32_47), .win4(wout32_48),
                    .aout1(aout33_48), .aout2(aout34_48), .aout3(aout35_48), .aout4(aout36_48),
                    .wout1(wout36_45), .wout2(wout36_46), .wout3(wout36_47), .wout4(wout36_48),
                    .sout11(sout33_45), .sout12(sout33_46), .sout13(sout33_47), .sout14(sout33_48),
                    .sout21(sout34_45), .sout22(sout34_46), .sout23(sout34_47), .sout24(sout34_48),
                    .sout31(sout35_45), .sout32(sout35_46), .sout33(sout35_47), .sout34(sout35_48),
                    .sout41(sout36_45), .sout42(sout36_46), .sout43(sout36_47), .sout44(sout36_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_9_13 (.clk(clk), .rst(rst),
                    .ain1(aout33_48), .ain2(aout34_48), .ain3(aout35_48), .ain4(aout36_48),
                    .win1(wout32_49), .win2(wout32_50), .win3(wout32_51), .win4(wout32_52),
                    .aout1(aout33_52), .aout2(aout34_52), .aout3(aout35_52), .aout4(aout36_52),
                    .wout1(wout36_49), .wout2(wout36_50), .wout3(wout36_51), .wout4(wout36_52),
                    .sout11(sout33_49), .sout12(sout33_50), .sout13(sout33_51), .sout14(sout33_52),
                    .sout21(sout34_49), .sout22(sout34_50), .sout23(sout34_51), .sout24(sout34_52),
                    .sout31(sout35_49), .sout32(sout35_50), .sout33(sout35_51), .sout34(sout35_52),
                    .sout41(sout36_49), .sout42(sout36_50), .sout43(sout36_51), .sout44(sout36_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_9_14 (.clk(clk), .rst(rst),
                    .ain1(aout33_52), .ain2(aout34_52), .ain3(aout35_52), .ain4(aout36_52),
                    .win1(wout32_53), .win2(wout32_54), .win3(wout32_55), .win4(wout32_56),
                    .aout1(aout33_56), .aout2(aout34_56), .aout3(aout35_56), .aout4(aout36_56),
                    .wout1(wout36_53), .wout2(wout36_54), .wout3(wout36_55), .wout4(wout36_56),
                    .sout11(sout33_53), .sout12(sout33_54), .sout13(sout33_55), .sout14(sout33_56),
                    .sout21(sout34_53), .sout22(sout34_54), .sout23(sout34_55), .sout24(sout34_56),
                    .sout31(sout35_53), .sout32(sout35_54), .sout33(sout35_55), .sout34(sout35_56),
                    .sout41(sout36_53), .sout42(sout36_54), .sout43(sout36_55), .sout44(sout36_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_9_15 (.clk(clk), .rst(rst),
                    .ain1(aout33_56), .ain2(aout34_56), .ain3(aout35_56), .ain4(aout36_56),
                    .win1(wout32_57), .win2(wout32_58), .win3(wout32_59), .win4(wout32_60),
                    .aout1(aout33_60), .aout2(aout34_60), .aout3(aout35_60), .aout4(aout36_60),
                    .wout1(wout36_57), .wout2(wout36_58), .wout3(wout36_59), .wout4(wout36_60),
                    .sout11(sout33_57), .sout12(sout33_58), .sout13(sout33_59), .sout14(sout33_60),
                    .sout21(sout34_57), .sout22(sout34_58), .sout23(sout34_59), .sout24(sout34_60),
                    .sout31(sout35_57), .sout32(sout35_58), .sout33(sout35_59), .sout34(sout35_60),
                    .sout41(sout36_57), .sout42(sout36_58), .sout43(sout36_59), .sout44(sout36_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_9_16 (.clk(clk), .rst(rst),
                    .ain1(aout33_60), .ain2(aout34_60), .ain3(aout35_60), .ain4(aout36_60),
                    .win1(wout32_61), .win2(wout32_62), .win3(wout32_63), .win4(wout32_64),
                    .aout1(aout33_64), .aout2(aout34_64), .aout3(aout35_64), .aout4(aout36_64),
                    .wout1(wout36_61), .wout2(wout36_62), .wout3(wout36_63), .wout4(wout36_64),
                    .sout11(sout33_61), .sout12(sout33_62), .sout13(sout33_63), .sout14(sout33_64),
                    .sout21(sout34_61), .sout22(sout34_62), .sout23(sout34_63), .sout24(sout34_64),
                    .sout31(sout35_61), .sout32(sout35_62), .sout33(sout35_63), .sout34(sout35_64),
                    .sout41(sout36_61), .sout42(sout36_62), .sout43(sout36_63), .sout44(sout36_64)
                    ); //4x4 MAC array
                    
                    
 
    //row10
    mac_array_4x4 mac_array_4x4_10_1 (.clk(clk), .rst(rst),
                    .ain1(ain37), .ain2(ain38), .ain3(ain39), .ain4(ain40),
                    .win1(wout36_1), .win2(wout36_2), .win3(wout36_3), .win4(wout36_4),
                    .aout1(aout37_4), .aout2(aout38_4), .aout3(aout39_4), .aout4(aout40_4),
                    .wout1(wout40_1), .wout2(wout40_2), .wout3(wout40_3), .wout4(wout40_4),
                    .sout11(sout37_1), .sout12(sout37_2), .sout13(sout37_3), .sout14(sout37_4),
                    .sout21(sout38_1), .sout22(sout38_2), .sout23(sout38_3), .sout24(sout38_4),
                    .sout31(sout39_1), .sout32(sout39_2), .sout33(sout39_3), .sout34(sout39_4),
                    .sout41(sout40_1), .sout42(sout40_2), .sout43(sout40_3), .sout44(sout40_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_10_2 (.clk(clk), .rst(rst),
                    .ain1(aout37_4), .ain2(aout38_4), .ain3(aout39_4), .ain4(aout40_4),
                    .win1(wout36_5), .win2(wout36_6), .win3(wout36_7), .win4(wout36_8),
                    .aout1(aout37_8), .aout2(aout38_8), .aout3(aout39_8), .aout4(aout40_8),
                    .wout1(wout40_5), .wout2(wout40_6), .wout3(wout40_7), .wout4(wout40_8),
                    .sout11(sout37_5), .sout12(sout37_6), .sout13(sout37_7), .sout14(sout37_8),
                    .sout21(sout38_5), .sout22(sout38_6), .sout23(sout38_7), .sout24(sout38_8),
                    .sout31(sout39_5), .sout32(sout39_6), .sout33(sout39_7), .sout34(sout39_8),
                    .sout41(sout40_5), .sout42(sout40_6), .sout43(sout40_7), .sout44(sout40_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_10_3 (.clk(clk), .rst(rst),
                    .ain1(aout37_8), .ain2(aout38_8), .ain3(aout39_8), .ain4(aout40_8),
                    .win1(wout36_9), .win2(wout36_10), .win3(wout36_11), .win4(wout36_12),
                    .aout1(aout37_12), .aout2(aout38_12), .aout3(aout39_12), .aout4(aout40_12),
                    .wout1(wout40_9), .wout2(wout40_10), .wout3(wout40_11), .wout4(wout40_12),
                    .sout11(sout37_9), .sout12(sout37_10), .sout13(sout37_11), .sout14(sout37_12),
                    .sout21(sout38_9), .sout22(sout38_10), .sout23(sout38_11), .sout24(sout38_12),
                    .sout31(sout39_9), .sout32(sout39_10), .sout33(sout39_11), .sout34(sout39_12),
                    .sout41(sout40_9), .sout42(sout40_10), .sout43(sout40_11), .sout44(sout40_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_10_4 (.clk(clk), .rst(rst),
                    .ain1(aout37_12), .ain2(aout38_12), .ain3(aout39_12), .ain4(aout40_12),
                    .win1(wout36_13), .win2(wout36_14), .win3(wout36_15), .win4(wout36_16),
                    .aout1(aout37_16), .aout2(aout38_16), .aout3(aout39_16), .aout4(aout40_16),
                    .wout1(wout40_13), .wout2(wout40_14), .wout3(wout40_15), .wout4(wout40_16),
                    .sout11(sout37_13), .sout12(sout37_14), .sout13(sout37_15), .sout14(sout37_16),
                    .sout21(sout38_13), .sout22(sout38_14), .sout23(sout38_15), .sout24(sout38_16),
                    .sout31(sout39_13), .sout32(sout39_14), .sout33(sout39_15), .sout34(sout39_16),
                    .sout41(sout40_13), .sout42(sout40_14), .sout43(sout40_15), .sout44(sout40_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_10_5 (.clk(clk), .rst(rst),
                    .ain1(aout37_16), .ain2(aout38_16), .ain3(aout39_16), .ain4(aout40_16),
                    .win1(wout36_17), .win2(wout36_18), .win3(wout36_19), .win4(wout36_20),
                    .aout1(aout37_20), .aout2(aout38_20), .aout3(aout39_20), .aout4(aout40_20),
                    .wout1(wout40_17), .wout2(wout40_18), .wout3(wout40_19), .wout4(wout40_20),
                    .sout11(sout37_17), .sout12(sout37_18), .sout13(sout37_19), .sout14(sout37_20),
                    .sout21(sout38_17), .sout22(sout38_18), .sout23(sout38_19), .sout24(sout38_20),
                    .sout31(sout39_17), .sout32(sout39_18), .sout33(sout39_19), .sout34(sout39_20),
                    .sout41(sout40_17), .sout42(sout40_18), .sout43(sout40_19), .sout44(sout40_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_10_6 (.clk(clk), .rst(rst),
                    .ain1(aout37_20), .ain2(aout38_20), .ain3(aout39_20), .ain4(aout40_20),
                    .win1(wout36_21), .win2(wout36_22), .win3(wout36_23), .win4(wout36_24),
                    .aout1(aout37_24), .aout2(aout38_24), .aout3(aout39_24), .aout4(aout40_24),
                    .wout1(wout40_21), .wout2(wout40_22), .wout3(wout40_23), .wout4(wout40_24),
                    .sout11(sout37_21), .sout12(sout37_22), .sout13(sout37_23), .sout14(sout37_24),
                    .sout21(sout38_21), .sout22(sout38_22), .sout23(sout38_23), .sout24(sout38_24),
                    .sout31(sout39_21), .sout32(sout39_22), .sout33(sout39_23), .sout34(sout39_24),
                    .sout41(sout40_21), .sout42(sout40_22), .sout43(sout40_23), .sout44(sout40_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_10_7 (.clk(clk), .rst(rst),
                    .ain1(aout37_24), .ain2(aout38_24), .ain3(aout39_24), .ain4(aout40_24),
                    .win1(wout36_25), .win2(wout36_26), .win3(wout36_27), .win4(wout36_28),
                    .aout1(aout37_28), .aout2(aout38_28), .aout3(aout39_28), .aout4(aout40_28),
                    .wout1(wout40_25), .wout2(wout40_26), .wout3(wout40_27), .wout4(wout40_28),
                    .sout11(sout37_25), .sout12(sout37_26), .sout13(sout37_27), .sout14(sout37_28),
                    .sout21(sout38_25), .sout22(sout38_26), .sout23(sout38_27), .sout24(sout38_28),
                    .sout31(sout39_25), .sout32(sout39_26), .sout33(sout39_27), .sout34(sout39_28),
                    .sout41(sout40_25), .sout42(sout40_26), .sout43(sout40_27), .sout44(sout40_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_10_8 (.clk(clk), .rst(rst),
                    .ain1(aout37_28), .ain2(aout38_28), .ain3(aout39_28), .ain4(aout40_28),
                    .win1(wout36_29), .win2(wout36_30), .win3(wout36_31), .win4(wout36_32),
                    .aout1(aout37_32), .aout2(aout38_32), .aout3(aout39_32), .aout4(aout40_32),
                    .wout1(wout40_29), .wout2(wout40_30), .wout3(wout40_31), .wout4(wout40_32),
                    .sout11(sout37_29), .sout12(sout37_30), .sout13(sout37_31), .sout14(sout37_32),
                    .sout21(sout38_29), .sout22(sout38_30), .sout23(sout38_31), .sout24(sout38_32),
                    .sout31(sout39_29), .sout32(sout39_30), .sout33(sout39_31), .sout34(sout39_32),
                    .sout41(sout40_29), .sout42(sout40_30), .sout43(sout40_31), .sout44(sout40_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_10_9 (.clk(clk), .rst(rst),
                    .ain1(aout37_32), .ain2(aout38_32), .ain3(aout39_32), .ain4(aout40_32),
                    .win1(wout36_33), .win2(wout36_34), .win3(wout36_35), .win4(wout36_36),
                    .aout1(aout37_36), .aout2(aout38_36), .aout3(aout39_36), .aout4(aout40_36),
                    .wout1(wout40_33), .wout2(wout40_34), .wout3(wout40_35), .wout4(wout40_36),
                    .sout11(sout37_33), .sout12(sout37_34), .sout13(sout37_35), .sout14(sout37_36),
                    .sout21(sout38_33), .sout22(sout38_34), .sout23(sout38_35), .sout24(sout38_36),
                    .sout31(sout39_33), .sout32(sout39_34), .sout33(sout39_35), .sout34(sout39_36),
                    .sout41(sout40_33), .sout42(sout40_34), .sout43(sout40_35), .sout44(sout40_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_10_10 (.clk(clk), .rst(rst),
                    .ain1(aout37_36), .ain2(aout38_36), .ain3(aout39_36), .ain4(aout40_36),
                    .win1(wout36_37), .win2(wout36_38), .win3(wout36_39), .win4(wout36_40),
                    .aout1(aout37_40), .aout2(aout38_40), .aout3(aout39_40), .aout4(aout40_40),
                    .wout1(wout40_37), .wout2(wout40_38), .wout3(wout40_39), .wout4(wout40_40),
                    .sout11(sout37_37), .sout12(sout37_38), .sout13(sout37_39), .sout14(sout37_40),
                    .sout21(sout38_37), .sout22(sout38_38), .sout23(sout38_39), .sout24(sout38_40),
                    .sout31(sout39_37), .sout32(sout39_38), .sout33(sout39_39), .sout34(sout39_40),
                    .sout41(sout40_37), .sout42(sout40_38), .sout43(sout40_39), .sout44(sout40_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_10_11 (.clk(clk), .rst(rst),
                    .ain1(aout37_40), .ain2(aout38_40), .ain3(aout39_40), .ain4(aout40_40),
                    .win1(wout36_41), .win2(wout36_42), .win3(wout36_43), .win4(wout36_44),
                    .aout1(aout37_44), .aout2(aout38_44), .aout3(aout39_44), .aout4(aout40_44),
                    .wout1(wout40_41), .wout2(wout40_42), .wout3(wout40_43), .wout4(wout40_44),
                    .sout11(sout37_41), .sout12(sout37_42), .sout13(sout37_43), .sout14(sout37_44),
                    .sout21(sout38_41), .sout22(sout38_42), .sout23(sout38_43), .sout24(sout38_44),
                    .sout31(sout39_41), .sout32(sout39_42), .sout33(sout39_43), .sout34(sout39_44),
                    .sout41(sout40_41), .sout42(sout40_42), .sout43(sout40_43), .sout44(sout40_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_10_12 (.clk(clk), .rst(rst),
                    .ain1(aout37_44), .ain2(aout38_44), .ain3(aout39_44), .ain4(aout40_44),
                    .win1(wout36_45), .win2(wout36_46), .win3(wout36_47), .win4(wout36_48),
                    .aout1(aout37_48), .aout2(aout38_48), .aout3(aout39_48), .aout4(aout40_48),
                    .wout1(wout40_45), .wout2(wout40_46), .wout3(wout40_47), .wout4(wout40_48),
                    .sout11(sout37_45), .sout12(sout37_46), .sout13(sout37_47), .sout14(sout37_48),
                    .sout21(sout38_45), .sout22(sout38_46), .sout23(sout38_47), .sout24(sout38_48),
                    .sout31(sout39_45), .sout32(sout39_46), .sout33(sout39_47), .sout34(sout39_48),
                    .sout41(sout40_45), .sout42(sout40_46), .sout43(sout40_47), .sout44(sout40_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_10_13 (.clk(clk), .rst(rst),
                    .ain1(aout37_48), .ain2(aout38_48), .ain3(aout39_48), .ain4(aout40_48),
                    .win1(wout36_49), .win2(wout36_50), .win3(wout36_51), .win4(wout36_52),
                    .aout1(aout37_52), .aout2(aout38_52), .aout3(aout39_52), .aout4(aout40_52),
                    .wout1(wout40_49), .wout2(wout40_50), .wout3(wout40_51), .wout4(wout40_52),
                    .sout11(sout37_49), .sout12(sout37_50), .sout13(sout37_51), .sout14(sout37_52),
                    .sout21(sout38_49), .sout22(sout38_50), .sout23(sout38_51), .sout24(sout38_52),
                    .sout31(sout39_49), .sout32(sout39_50), .sout33(sout39_51), .sout34(sout39_52),
                    .sout41(sout40_49), .sout42(sout40_50), .sout43(sout40_51), .sout44(sout40_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_10_14 (.clk(clk), .rst(rst),
                    .ain1(aout37_52), .ain2(aout38_52), .ain3(aout39_52), .ain4(aout40_52),
                    .win1(wout36_53), .win2(wout36_54), .win3(wout36_55), .win4(wout36_56),
                    .aout1(aout37_56), .aout2(aout38_56), .aout3(aout39_56), .aout4(aout40_56),
                    .wout1(wout40_53), .wout2(wout40_54), .wout3(wout40_55), .wout4(wout40_56),
                    .sout11(sout37_53), .sout12(sout37_54), .sout13(sout37_55), .sout14(sout37_56),
                    .sout21(sout38_53), .sout22(sout38_54), .sout23(sout38_55), .sout24(sout38_56),
                    .sout31(sout39_53), .sout32(sout39_54), .sout33(sout39_55), .sout34(sout39_56),
                    .sout41(sout40_53), .sout42(sout40_54), .sout43(sout40_55), .sout44(sout40_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_10_15 (.clk(clk), .rst(rst),
                    .ain1(aout37_56), .ain2(aout38_56), .ain3(aout39_56), .ain4(aout40_56),
                    .win1(wout36_57), .win2(wout36_58), .win3(wout36_59), .win4(wout36_60),
                    .aout1(aout37_60), .aout2(aout38_60), .aout3(aout39_60), .aout4(aout40_60),
                    .wout1(wout40_57), .wout2(wout40_58), .wout3(wout40_59), .wout4(wout40_60),
                    .sout11(sout37_57), .sout12(sout37_58), .sout13(sout37_59), .sout14(sout37_60),
                    .sout21(sout38_57), .sout22(sout38_58), .sout23(sout38_59), .sout24(sout38_60),
                    .sout31(sout39_57), .sout32(sout39_58), .sout33(sout39_59), .sout34(sout39_60),
                    .sout41(sout40_57), .sout42(sout40_58), .sout43(sout40_59), .sout44(sout40_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_10_16 (.clk(clk), .rst(rst),
                    .ain1(aout37_60), .ain2(aout38_60), .ain3(aout39_60), .ain4(aout40_60),
                    .win1(wout36_61), .win2(wout36_62), .win3(wout36_63), .win4(wout36_64),
                    .aout1(aout37_64), .aout2(aout38_64), .aout3(aout39_64), .aout4(aout40_64),
                    .wout1(wout40_61), .wout2(wout40_62), .wout3(wout40_63), .wout4(wout40_64),
                    .sout11(sout37_61), .sout12(sout37_62), .sout13(sout37_63), .sout14(sout37_64),
                    .sout21(sout38_61), .sout22(sout38_62), .sout23(sout38_63), .sout24(sout38_64),
                    .sout31(sout39_61), .sout32(sout39_62), .sout33(sout39_63), .sout34(sout39_64),
                    .sout41(sout40_61), .sout42(sout40_62), .sout43(sout40_63), .sout44(sout40_64)
                    ); //4x4 MAC array
                    
                 
    //row11
    mac_array_4x4 mac_array_4x4_11_1 (.clk(clk), .rst(rst),
                    .ain1(ain41), .ain2(ain42), .ain3(ain43), .ain4(ain44),
                    .win1(wout40_1), .win2(wout40_2), .win3(wout40_3), .win4(wout40_4),
                    .aout1(aout41_4), .aout2(aout42_4), .aout3(aout43_4), .aout4(aout44_4),
                    .wout1(wout44_1), .wout2(wout44_2), .wout3(wout44_3), .wout4(wout44_4),
                    .sout11(sout41_1), .sout12(sout41_2), .sout13(sout41_3), .sout14(sout41_4),
                    .sout21(sout42_1), .sout22(sout42_2), .sout23(sout42_3), .sout24(sout42_4),
                    .sout31(sout43_1), .sout32(sout43_2), .sout33(sout43_3), .sout34(sout43_4),
                    .sout41(sout44_1), .sout42(sout44_2), .sout43(sout44_3), .sout44(sout44_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_11_2 (.clk(clk), .rst(rst),
                    .ain1(aout41_4), .ain2(aout42_4), .ain3(aout43_4), .ain4(aout44_4),
                    .win1(wout40_5), .win2(wout40_6), .win3(wout40_7), .win4(wout40_8),
                    .aout1(aout41_8), .aout2(aout42_8), .aout3(aout43_8), .aout4(aout44_8),
                    .wout1(wout44_5), .wout2(wout44_6), .wout3(wout44_7), .wout4(wout44_8),
                    .sout11(sout41_5), .sout12(sout41_6), .sout13(sout41_7), .sout14(sout41_8),
                    .sout21(sout42_5), .sout22(sout42_6), .sout23(sout42_7), .sout24(sout42_8),
                    .sout31(sout43_5), .sout32(sout43_6), .sout33(sout43_7), .sout34(sout43_8),
                    .sout41(sout44_5), .sout42(sout44_6), .sout43(sout44_7), .sout44(sout44_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_11_3 (.clk(clk), .rst(rst),
                    .ain1(aout41_8), .ain2(aout42_8), .ain3(aout43_8), .ain4(aout44_8),
                    .win1(wout40_9), .win2(wout40_10), .win3(wout40_11), .win4(wout40_12),
                    .aout1(aout41_12), .aout2(aout42_12), .aout3(aout43_12), .aout4(aout44_12),
                    .wout1(wout44_9), .wout2(wout44_10), .wout3(wout44_11), .wout4(wout44_12),
                    .sout11(sout41_9), .sout12(sout41_10), .sout13(sout41_11), .sout14(sout41_12),
                    .sout21(sout42_9), .sout22(sout42_10), .sout23(sout42_11), .sout24(sout42_12),
                    .sout31(sout43_9), .sout32(sout43_10), .sout33(sout43_11), .sout34(sout43_12),
                    .sout41(sout44_9), .sout42(sout44_10), .sout43(sout44_11), .sout44(sout44_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_11_4 (.clk(clk), .rst(rst),
                    .ain1(aout41_12), .ain2(aout42_12), .ain3(aout43_12), .ain4(aout44_12),
                    .win1(wout40_13), .win2(wout40_14), .win3(wout40_15), .win4(wout40_16),
                    .aout1(aout41_16), .aout2(aout42_16), .aout3(aout43_16), .aout4(aout44_16),
                    .wout1(wout44_13), .wout2(wout44_14), .wout3(wout44_15), .wout4(wout44_16),
                    .sout11(sout41_13), .sout12(sout41_14), .sout13(sout41_15), .sout14(sout41_16),
                    .sout21(sout42_13), .sout22(sout42_14), .sout23(sout42_15), .sout24(sout42_16),
                    .sout31(sout43_13), .sout32(sout43_14), .sout33(sout43_15), .sout34(sout43_16),
                    .sout41(sout44_13), .sout42(sout44_14), .sout43(sout44_15), .sout44(sout44_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_11_5 (.clk(clk), .rst(rst),
                    .ain1(aout41_16), .ain2(aout42_16), .ain3(aout43_16), .ain4(aout44_16),
                    .win1(wout40_17), .win2(wout40_18), .win3(wout40_19), .win4(wout40_20),
                    .aout1(aout41_20), .aout2(aout42_20), .aout3(aout43_20), .aout4(aout44_20),
                    .wout1(wout44_17), .wout2(wout44_18), .wout3(wout44_19), .wout4(wout44_20),
                    .sout11(sout41_17), .sout12(sout41_18), .sout13(sout41_19), .sout14(sout41_20),
                    .sout21(sout42_17), .sout22(sout42_18), .sout23(sout42_19), .sout24(sout42_20),
                    .sout31(sout43_17), .sout32(sout43_18), .sout33(sout43_19), .sout34(sout43_20),
                    .sout41(sout44_17), .sout42(sout44_18), .sout43(sout44_19), .sout44(sout44_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_11_6 (.clk(clk), .rst(rst),
                    .ain1(aout41_20), .ain2(aout42_20), .ain3(aout43_20), .ain4(aout44_20),
                    .win1(wout40_21), .win2(wout40_22), .win3(wout40_23), .win4(wout40_24),
                    .aout1(aout41_24), .aout2(aout42_24), .aout3(aout43_24), .aout4(aout44_24),
                    .wout1(wout44_21), .wout2(wout44_22), .wout3(wout44_23), .wout4(wout44_24),
                    .sout11(sout41_21), .sout12(sout41_22), .sout13(sout41_23), .sout14(sout41_24),
                    .sout21(sout42_21), .sout22(sout42_22), .sout23(sout42_23), .sout24(sout42_24),
                    .sout31(sout43_21), .sout32(sout43_22), .sout33(sout43_23), .sout34(sout43_24),
                    .sout41(sout44_21), .sout42(sout44_22), .sout43(sout44_23), .sout44(sout44_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_11_7 (.clk(clk), .rst(rst),
                    .ain1(aout41_24), .ain2(aout42_24), .ain3(aout43_24), .ain4(aout44_24),
                    .win1(wout40_25), .win2(wout40_26), .win3(wout40_27), .win4(wout40_28),
                    .aout1(aout41_28), .aout2(aout42_28), .aout3(aout43_28), .aout4(aout44_28),
                    .wout1(wout44_25), .wout2(wout44_26), .wout3(wout44_27), .wout4(wout44_28),
                    .sout11(sout41_25), .sout12(sout41_26), .sout13(sout41_27), .sout14(sout41_28),
                    .sout21(sout42_25), .sout22(sout42_26), .sout23(sout42_27), .sout24(sout42_28),
                    .sout31(sout43_25), .sout32(sout43_26), .sout33(sout43_27), .sout34(sout43_28),
                    .sout41(sout44_25), .sout42(sout44_26), .sout43(sout44_27), .sout44(sout44_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_11_8 (.clk(clk), .rst(rst),
                    .ain1(aout41_28), .ain2(aout42_28), .ain3(aout43_28), .ain4(aout44_28),
                    .win1(wout40_29), .win2(wout40_30), .win3(wout40_31), .win4(wout40_32),
                    .aout1(aout41_32), .aout2(aout42_32), .aout3(aout43_32), .aout4(aout44_32),
                    .wout1(wout44_29), .wout2(wout44_30), .wout3(wout44_31), .wout4(wout44_32),
                    .sout11(sout41_29), .sout12(sout41_30), .sout13(sout41_31), .sout14(sout41_32),
                    .sout21(sout42_29), .sout22(sout42_30), .sout23(sout42_31), .sout24(sout42_32),
                    .sout31(sout43_29), .sout32(sout43_30), .sout33(sout43_31), .sout34(sout43_32),
                    .sout41(sout44_29), .sout42(sout44_30), .sout43(sout44_31), .sout44(sout44_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_11_9 (.clk(clk), .rst(rst),
                    .ain1(aout41_32), .ain2(aout42_32), .ain3(aout43_32), .ain4(aout44_32),
                    .win1(wout40_33), .win2(wout40_34), .win3(wout40_35), .win4(wout40_36),
                    .aout1(aout41_36), .aout2(aout42_36), .aout3(aout43_36), .aout4(aout44_36),
                    .wout1(wout44_33), .wout2(wout44_34), .wout3(wout44_35), .wout4(wout44_36),
                    .sout11(sout41_33), .sout12(sout41_34), .sout13(sout41_35), .sout14(sout41_36),
                    .sout21(sout42_33), .sout22(sout42_34), .sout23(sout42_35), .sout24(sout42_36),
                    .sout31(sout43_33), .sout32(sout43_34), .sout33(sout43_35), .sout34(sout43_36),
                    .sout41(sout44_33), .sout42(sout44_34), .sout43(sout44_35), .sout44(sout44_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_11_10 (.clk(clk), .rst(rst),
                    .ain1(aout41_36), .ain2(aout42_36), .ain3(aout43_36), .ain4(aout44_36),
                    .win1(wout40_37), .win2(wout40_38), .win3(wout40_39), .win4(wout40_40),
                    .aout1(aout41_40), .aout2(aout42_40), .aout3(aout43_40), .aout4(aout44_40),
                    .wout1(wout44_37), .wout2(wout44_38), .wout3(wout44_39), .wout4(wout44_40),
                    .sout11(sout41_37), .sout12(sout41_38), .sout13(sout41_39), .sout14(sout41_40),
                    .sout21(sout42_37), .sout22(sout42_38), .sout23(sout42_39), .sout24(sout42_40),
                    .sout31(sout43_37), .sout32(sout43_38), .sout33(sout43_39), .sout34(sout43_40),
                    .sout41(sout44_37), .sout42(sout44_38), .sout43(sout44_39), .sout44(sout44_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_11_11 (.clk(clk), .rst(rst),
                    .ain1(aout41_40), .ain2(aout42_40), .ain3(aout43_40), .ain4(aout44_40),
                    .win1(wout40_41), .win2(wout40_42), .win3(wout40_43), .win4(wout40_44),
                    .aout1(aout41_44), .aout2(aout42_44), .aout3(aout43_44), .aout4(aout44_44),
                    .wout1(wout44_41), .wout2(wout44_42), .wout3(wout44_43), .wout4(wout44_44),
                    .sout11(sout41_41), .sout12(sout41_42), .sout13(sout41_43), .sout14(sout41_44),
                    .sout21(sout42_41), .sout22(sout42_42), .sout23(sout42_43), .sout24(sout42_44),
                    .sout31(sout43_41), .sout32(sout43_42), .sout33(sout43_43), .sout34(sout43_44),
                    .sout41(sout44_41), .sout42(sout44_42), .sout43(sout44_43), .sout44(sout44_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_11_12 (.clk(clk), .rst(rst),
                    .ain1(aout41_44), .ain2(aout42_44), .ain3(aout43_44), .ain4(aout44_44),
                    .win1(wout40_45), .win2(wout40_46), .win3(wout40_47), .win4(wout40_48),
                    .aout1(aout41_48), .aout2(aout42_48), .aout3(aout43_48), .aout4(aout44_48),
                    .wout1(wout44_45), .wout2(wout44_46), .wout3(wout44_47), .wout4(wout44_48),
                    .sout11(sout41_45), .sout12(sout41_46), .sout13(sout41_47), .sout14(sout41_48),
                    .sout21(sout42_45), .sout22(sout42_46), .sout23(sout42_47), .sout24(sout42_48),
                    .sout31(sout43_45), .sout32(sout43_46), .sout33(sout43_47), .sout34(sout43_48),
                    .sout41(sout44_45), .sout42(sout44_46), .sout43(sout44_47), .sout44(sout44_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_11_13 (.clk(clk), .rst(rst),
                    .ain1(aout41_48), .ain2(aout42_48), .ain3(aout43_48), .ain4(aout44_48),
                    .win1(wout40_49), .win2(wout40_50), .win3(wout40_51), .win4(wout40_52),
                    .aout1(aout41_52), .aout2(aout42_52), .aout3(aout43_52), .aout4(aout44_52),
                    .wout1(wout44_49), .wout2(wout44_50), .wout3(wout44_51), .wout4(wout44_52),
                    .sout11(sout41_49), .sout12(sout41_50), .sout13(sout41_51), .sout14(sout41_52),
                    .sout21(sout42_49), .sout22(sout42_50), .sout23(sout42_51), .sout24(sout42_52),
                    .sout31(sout43_49), .sout32(sout43_50), .sout33(sout43_51), .sout34(sout43_52),
                    .sout41(sout44_49), .sout42(sout44_50), .sout43(sout44_51), .sout44(sout44_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_11_14 (.clk(clk), .rst(rst),
                    .ain1(aout41_52), .ain2(aout42_52), .ain3(aout43_52), .ain4(aout44_52),
                    .win1(wout40_53), .win2(wout40_54), .win3(wout40_55), .win4(wout40_56),
                    .aout1(aout41_56), .aout2(aout42_56), .aout3(aout43_56), .aout4(aout44_56),
                    .wout1(wout44_53), .wout2(wout44_54), .wout3(wout44_55), .wout4(wout44_56),
                    .sout11(sout41_53), .sout12(sout41_54), .sout13(sout41_55), .sout14(sout41_56),
                    .sout21(sout42_53), .sout22(sout42_54), .sout23(sout42_55), .sout24(sout42_56),
                    .sout31(sout43_53), .sout32(sout43_54), .sout33(sout43_55), .sout34(sout43_56),
                    .sout41(sout44_53), .sout42(sout44_54), .sout43(sout44_55), .sout44(sout44_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_11_15 (.clk(clk), .rst(rst),
                    .ain1(aout41_56), .ain2(aout42_56), .ain3(aout43_56), .ain4(aout44_56),
                    .win1(wout40_57), .win2(wout40_58), .win3(wout40_59), .win4(wout40_60),
                    .aout1(aout41_60), .aout2(aout42_60), .aout3(aout43_60), .aout4(aout44_60),
                    .wout1(wout44_57), .wout2(wout44_58), .wout3(wout44_59), .wout4(wout44_60),
                    .sout11(sout41_57), .sout12(sout41_58), .sout13(sout41_59), .sout14(sout41_60),
                    .sout21(sout42_57), .sout22(sout42_58), .sout23(sout42_59), .sout24(sout42_60),
                    .sout31(sout43_57), .sout32(sout43_58), .sout33(sout43_59), .sout34(sout43_60),
                    .sout41(sout44_57), .sout42(sout44_58), .sout43(sout44_59), .sout44(sout44_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_11_16 (.clk(clk), .rst(rst),
                    .ain1(aout41_60), .ain2(aout42_60), .ain3(aout43_60), .ain4(aout44_60),
                    .win1(wout40_61), .win2(wout40_62), .win3(wout40_63), .win4(wout40_64),
                    .aout1(aout41_64), .aout2(aout42_64), .aout3(aout43_64), .aout4(aout44_64),
                    .wout1(wout44_61), .wout2(wout44_62), .wout3(wout44_63), .wout4(wout44_64),
                    .sout11(sout41_61), .sout12(sout41_62), .sout13(sout41_63), .sout14(sout41_64),
                    .sout21(sout42_61), .sout22(sout42_62), .sout23(sout42_63), .sout24(sout42_64),
                    .sout31(sout43_61), .sout32(sout43_62), .sout33(sout43_63), .sout34(sout43_64),
                    .sout41(sout44_61), .sout42(sout44_62), .sout43(sout44_63), .sout44(sout44_64)
                    ); //4x4 MAC array
                    
              
    mac_array_4x4 mac_array_4x4_12_1 (.clk(clk), .rst(rst),
                    .ain1(ain45), .ain2(ain46), .ain3(ain47), .ain4(ain48),
                    .win1(wout44_1), .win2(wout44_2), .win3(wout44_3), .win4(wout44_4),
                    .aout1(aout45_4), .aout2(aout46_4), .aout3(aout47_4), .aout4(aout48_4),
                    .wout1(wout48_1), .wout2(wout48_2), .wout3(wout48_3), .wout4(wout48_4),
                    .sout11(sout45_1), .sout12(sout45_2), .sout13(sout45_3), .sout14(sout45_4),
                    .sout21(sout46_1), .sout22(sout46_2), .sout23(sout46_3), .sout24(sout46_4),
                    .sout31(sout47_1), .sout32(sout47_2), .sout33(sout47_3), .sout34(sout47_4),
                    .sout41(sout48_1), .sout42(sout48_2), .sout43(sout48_3), .sout44(sout48_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_12_2 (.clk(clk), .rst(rst),
                    .ain1(aout45_4), .ain2(aout46_4), .ain3(aout47_4), .ain4(aout48_4),
                    .win1(wout44_5), .win2(wout44_6), .win3(wout44_7), .win4(wout44_8),
                    .aout1(aout45_8), .aout2(aout46_8), .aout3(aout47_8), .aout4(aout48_8),
                    .wout1(wout48_5), .wout2(wout48_6), .wout3(wout48_7), .wout4(wout48_8),
                    .sout11(sout45_5), .sout12(sout45_6), .sout13(sout45_7), .sout14(sout45_8),
                    .sout21(sout46_5), .sout22(sout46_6), .sout23(sout46_7), .sout24(sout46_8),
                    .sout31(sout47_5), .sout32(sout47_6), .sout33(sout47_7), .sout34(sout47_8),
                    .sout41(sout48_5), .sout42(sout48_6), .sout43(sout48_7), .sout44(sout48_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_12_3 (.clk(clk), .rst(rst),
                    .ain1(aout45_8), .ain2(aout46_8), .ain3(aout47_8), .ain4(aout48_8),
                    .win1(wout44_9), .win2(wout44_10), .win3(wout44_11), .win4(wout44_12),
                    .aout1(aout45_12), .aout2(aout46_12), .aout3(aout47_12), .aout4(aout48_12),
                    .wout1(wout48_9), .wout2(wout48_10), .wout3(wout48_11), .wout4(wout48_12),
                    .sout11(sout45_9), .sout12(sout45_10), .sout13(sout45_11), .sout14(sout45_12),
                    .sout21(sout46_9), .sout22(sout46_10), .sout23(sout46_11), .sout24(sout46_12),
                    .sout31(sout47_9), .sout32(sout47_10), .sout33(sout47_11), .sout34(sout47_12),
                    .sout41(sout48_9), .sout42(sout48_10), .sout43(sout48_11), .sout44(sout48_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_12_4 (.clk(clk), .rst(rst),
                    .ain1(aout45_12), .ain2(aout46_12), .ain3(aout47_12), .ain4(aout48_12),
                    .win1(wout44_13), .win2(wout44_14), .win3(wout44_15), .win4(wout44_16),
                    .aout1(aout45_16), .aout2(aout46_16), .aout3(aout47_16), .aout4(aout48_16),
                    .wout1(wout48_13), .wout2(wout48_14), .wout3(wout48_15), .wout4(wout48_16),
                    .sout11(sout45_13), .sout12(sout45_14), .sout13(sout45_15), .sout14(sout45_16),
                    .sout21(sout46_13), .sout22(sout46_14), .sout23(sout46_15), .sout24(sout46_16),
                    .sout31(sout47_13), .sout32(sout47_14), .sout33(sout47_15), .sout34(sout47_16),
                    .sout41(sout48_13), .sout42(sout48_14), .sout43(sout48_15), .sout44(sout48_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_12_5 (.clk(clk), .rst(rst),
                    .ain1(aout45_16), .ain2(aout46_16), .ain3(aout47_16), .ain4(aout48_16),
                    .win1(wout44_17), .win2(wout44_18), .win3(wout44_19), .win4(wout44_20),
                    .aout1(aout45_20), .aout2(aout46_20), .aout3(aout47_20), .aout4(aout48_20),
                    .wout1(wout48_17), .wout2(wout48_18), .wout3(wout48_19), .wout4(wout48_20),
                    .sout11(sout45_17), .sout12(sout45_18), .sout13(sout45_19), .sout14(sout45_20),
                    .sout21(sout46_17), .sout22(sout46_18), .sout23(sout46_19), .sout24(sout46_20),
                    .sout31(sout47_17), .sout32(sout47_18), .sout33(sout47_19), .sout34(sout47_20),
                    .sout41(sout48_17), .sout42(sout48_18), .sout43(sout48_19), .sout44(sout48_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_12_6 (.clk(clk), .rst(rst),
                    .ain1(aout45_20), .ain2(aout46_20), .ain3(aout47_20), .ain4(aout48_20),
                    .win1(wout44_21), .win2(wout44_22), .win3(wout44_23), .win4(wout44_24),
                    .aout1(aout45_24), .aout2(aout46_24), .aout3(aout47_24), .aout4(aout48_24),
                    .wout1(wout48_21), .wout2(wout48_22), .wout3(wout48_23), .wout4(wout48_24),
                    .sout11(sout45_21), .sout12(sout45_22), .sout13(sout45_23), .sout14(sout45_24),
                    .sout21(sout46_21), .sout22(sout46_22), .sout23(sout46_23), .sout24(sout46_24),
                    .sout31(sout47_21), .sout32(sout47_22), .sout33(sout47_23), .sout34(sout47_24),
                    .sout41(sout48_21), .sout42(sout48_22), .sout43(sout48_23), .sout44(sout48_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_12_7 (.clk(clk), .rst(rst),
                    .ain1(aout45_24), .ain2(aout46_24), .ain3(aout47_24), .ain4(aout48_24),
                    .win1(wout44_25), .win2(wout44_26), .win3(wout44_27), .win4(wout44_28),
                    .aout1(aout45_28), .aout2(aout46_28), .aout3(aout47_28), .aout4(aout48_28),
                    .wout1(wout48_25), .wout2(wout48_26), .wout3(wout48_27), .wout4(wout48_28),
                    .sout11(sout45_25), .sout12(sout45_26), .sout13(sout45_27), .sout14(sout45_28),
                    .sout21(sout46_25), .sout22(sout46_26), .sout23(sout46_27), .sout24(sout46_28),
                    .sout31(sout47_25), .sout32(sout47_26), .sout33(sout47_27), .sout34(sout47_28),
                    .sout41(sout48_25), .sout42(sout48_26), .sout43(sout48_27), .sout44(sout48_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_12_8 (.clk(clk), .rst(rst),
                    .ain1(aout45_28), .ain2(aout46_28), .ain3(aout47_28), .ain4(aout48_28),
                    .win1(wout44_29), .win2(wout44_30), .win3(wout44_31), .win4(wout44_32),
                    .aout1(aout45_32), .aout2(aout46_32), .aout3(aout47_32), .aout4(aout48_32),
                    .wout1(wout48_29), .wout2(wout48_30), .wout3(wout48_31), .wout4(wout48_32),
                    .sout11(sout45_29), .sout12(sout45_30), .sout13(sout45_31), .sout14(sout45_32),
                    .sout21(sout46_29), .sout22(sout46_30), .sout23(sout46_31), .sout24(sout46_32),
                    .sout31(sout47_29), .sout32(sout47_30), .sout33(sout47_31), .sout34(sout47_32),
                    .sout41(sout48_29), .sout42(sout48_30), .sout43(sout48_31), .sout44(sout48_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_12_9 (.clk(clk), .rst(rst),
                    .ain1(aout45_32), .ain2(aout46_32), .ain3(aout47_32), .ain4(aout48_32),
                    .win1(wout44_33), .win2(wout44_34), .win3(wout44_35), .win4(wout44_36),
                    .aout1(aout45_36), .aout2(aout46_36), .aout3(aout47_36), .aout4(aout48_36),
                    .wout1(wout48_33), .wout2(wout48_34), .wout3(wout48_35), .wout4(wout48_36),
                    .sout11(sout45_33), .sout12(sout45_34), .sout13(sout45_35), .sout14(sout45_36),
                    .sout21(sout46_33), .sout22(sout46_34), .sout23(sout46_35), .sout24(sout46_36),
                    .sout31(sout47_33), .sout32(sout47_34), .sout33(sout47_35), .sout34(sout47_36),
                    .sout41(sout48_33), .sout42(sout48_34), .sout43(sout48_35), .sout44(sout48_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_12_10 (.clk(clk), .rst(rst),
                    .ain1(aout45_36), .ain2(aout46_36), .ain3(aout47_36), .ain4(aout48_36),
                    .win1(wout44_37), .win2(wout44_38), .win3(wout44_39), .win4(wout44_40),
                    .aout1(aout45_40), .aout2(aout46_40), .aout3(aout47_40), .aout4(aout48_40),
                    .wout1(wout48_37), .wout2(wout48_38), .wout3(wout48_39), .wout4(wout48_40),
                    .sout11(sout45_37), .sout12(sout45_38), .sout13(sout45_39), .sout14(sout45_40),
                    .sout21(sout46_37), .sout22(sout46_38), .sout23(sout46_39), .sout24(sout46_40),
                    .sout31(sout47_37), .sout32(sout47_38), .sout33(sout47_39), .sout34(sout47_40),
                    .sout41(sout48_37), .sout42(sout48_38), .sout43(sout48_39), .sout44(sout48_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_12_11 (.clk(clk), .rst(rst),
                    .ain1(aout45_40), .ain2(aout46_40), .ain3(aout47_40), .ain4(aout48_40),
                    .win1(wout44_41), .win2(wout44_42), .win3(wout44_43), .win4(wout44_44),
                    .aout1(aout45_44), .aout2(aout46_44), .aout3(aout47_44), .aout4(aout48_44),
                    .wout1(wout48_41), .wout2(wout48_42), .wout3(wout48_43), .wout4(wout48_44),
                    .sout11(sout45_41), .sout12(sout45_42), .sout13(sout45_43), .sout14(sout45_44),
                    .sout21(sout46_41), .sout22(sout46_42), .sout23(sout46_43), .sout24(sout46_44),
                    .sout31(sout47_41), .sout32(sout47_42), .sout33(sout47_43), .sout34(sout47_44),
                    .sout41(sout48_41), .sout42(sout48_42), .sout43(sout48_43), .sout44(sout48_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_12_12 (.clk(clk), .rst(rst),
                    .ain1(aout45_44), .ain2(aout46_44), .ain3(aout47_44), .ain4(aout48_44),
                    .win1(wout44_45), .win2(wout44_46), .win3(wout44_47), .win4(wout44_48),
                    .aout1(aout45_48), .aout2(aout46_48), .aout3(aout47_48), .aout4(aout48_48),
                    .wout1(wout48_45), .wout2(wout48_46), .wout3(wout48_47), .wout4(wout48_48),
                    .sout11(sout45_45), .sout12(sout45_46), .sout13(sout45_47), .sout14(sout45_48),
                    .sout21(sout46_45), .sout22(sout46_46), .sout23(sout46_47), .sout24(sout46_48),
                    .sout31(sout47_45), .sout32(sout47_46), .sout33(sout47_47), .sout34(sout47_48),
                    .sout41(sout48_45), .sout42(sout48_46), .sout43(sout48_47), .sout44(sout48_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_12_13 (.clk(clk), .rst(rst),
                    .ain1(aout45_48), .ain2(aout46_48), .ain3(aout47_48), .ain4(aout48_48),
                    .win1(wout44_49), .win2(wout44_50), .win3(wout44_51), .win4(wout44_52),
                    .aout1(aout45_52), .aout2(aout46_52), .aout3(aout47_52), .aout4(aout48_52),
                    .wout1(wout48_49), .wout2(wout48_50), .wout3(wout48_51), .wout4(wout48_52),
                    .sout11(sout45_49), .sout12(sout45_50), .sout13(sout45_51), .sout14(sout45_52),
                    .sout21(sout46_49), .sout22(sout46_50), .sout23(sout46_51), .sout24(sout46_52),
                    .sout31(sout47_49), .sout32(sout47_50), .sout33(sout47_51), .sout34(sout47_52),
                    .sout41(sout48_49), .sout42(sout48_50), .sout43(sout48_51), .sout44(sout48_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_12_14 (.clk(clk), .rst(rst),
                    .ain1(aout45_52), .ain2(aout46_52), .ain3(aout47_52), .ain4(aout48_52),
                    .win1(wout44_53), .win2(wout44_54), .win3(wout44_55), .win4(wout44_56),
                    .aout1(aout45_56), .aout2(aout46_56), .aout3(aout47_56), .aout4(aout48_56),
                    .wout1(wout48_53), .wout2(wout48_54), .wout3(wout48_55), .wout4(wout48_56),
                    .sout11(sout45_53), .sout12(sout45_54), .sout13(sout45_55), .sout14(sout45_56),
                    .sout21(sout46_53), .sout22(sout46_54), .sout23(sout46_55), .sout24(sout46_56),
                    .sout31(sout47_53), .sout32(sout47_54), .sout33(sout47_55), .sout34(sout47_56),
                    .sout41(sout48_53), .sout42(sout48_54), .sout43(sout48_55), .sout44(sout48_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_12_15 (.clk(clk), .rst(rst),
                    .ain1(aout45_56), .ain2(aout46_56), .ain3(aout47_56), .ain4(aout48_56),
                    .win1(wout44_57), .win2(wout44_58), .win3(wout44_59), .win4(wout44_60),
                    .aout1(aout45_60), .aout2(aout46_60), .aout3(aout47_60), .aout4(aout48_60),
                    .wout1(wout48_57), .wout2(wout48_58), .wout3(wout48_59), .wout4(wout48_60),
                    .sout11(sout45_57), .sout12(sout45_58), .sout13(sout45_59), .sout14(sout45_60),
                    .sout21(sout46_57), .sout22(sout46_58), .sout23(sout46_59), .sout24(sout46_60),
                    .sout31(sout47_57), .sout32(sout47_58), .sout33(sout47_59), .sout34(sout47_60),
                    .sout41(sout48_57), .sout42(sout48_58), .sout43(sout48_59), .sout44(sout48_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_12_16 (.clk(clk), .rst(rst),
                    .ain1(aout45_60), .ain2(aout46_60), .ain3(aout47_60), .ain4(aout48_60),
                    .win1(wout44_61), .win2(wout44_62), .win3(wout44_63), .win4(wout44_64),
                    .aout1(aout45_64), .aout2(aout46_64), .aout3(aout47_64), .aout4(aout48_64),
                    .wout1(wout48_61), .wout2(wout48_62), .wout3(wout48_63), .wout4(wout48_64),
                    .sout11(sout45_61), .sout12(sout45_62), .sout13(sout45_63), .sout14(sout45_64),
                    .sout21(sout46_61), .sout22(sout46_62), .sout23(sout46_63), .sout24(sout46_64),
                    .sout31(sout47_61), .sout32(sout47_62), .sout33(sout47_63), .sout34(sout47_64),
                    .sout41(sout48_61), .sout42(sout48_62), .sout43(sout48_63), .sout44(sout48_64)
                    ); //4x4 MAC array
                        
                            
                        
    //row13
    mac_array_4x4 mac_array_4x4_13_1 (.clk(clk), .rst(rst),
                    .ain1(ain49), .ain2(ain50), .ain3(ain51), .ain4(ain52),
                    .win1(wout48_1), .win2(wout48_2), .win3(wout48_3), .win4(wout48_4),
                    .aout1(aout49_4), .aout2(aout50_4), .aout3(aout51_4), .aout4(aout52_4),
                    .wout1(wout52_1), .wout2(wout52_2), .wout3(wout52_3), .wout4(wout52_4),
                    .sout11(sout49_1), .sout12(sout49_2), .sout13(sout49_3), .sout14(sout49_4),
                    .sout21(sout50_1), .sout22(sout50_2), .sout23(sout50_3), .sout24(sout50_4),
                    .sout31(sout51_1), .sout32(sout51_2), .sout33(sout51_3), .sout34(sout51_4),
                    .sout41(sout52_1), .sout42(sout52_2), .sout43(sout52_3), .sout44(sout52_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_13_2 (.clk(clk), .rst(rst),
                    .ain1(aout49_4), .ain2(aout50_4), .ain3(aout51_4), .ain4(aout52_4),
                    .win1(wout48_5), .win2(wout48_6), .win3(wout48_7), .win4(wout48_8),
                    .aout1(aout49_8), .aout2(aout50_8), .aout3(aout51_8), .aout4(aout52_8),
                    .wout1(wout52_5), .wout2(wout52_6), .wout3(wout52_7), .wout4(wout52_8),
                    .sout11(sout49_5), .sout12(sout49_6), .sout13(sout49_7), .sout14(sout49_8),
                    .sout21(sout50_5), .sout22(sout50_6), .sout23(sout50_7), .sout24(sout50_8),
                    .sout31(sout51_5), .sout32(sout51_6), .sout33(sout51_7), .sout34(sout51_8),
                    .sout41(sout52_5), .sout42(sout52_6), .sout43(sout52_7), .sout44(sout52_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_13_3 (.clk(clk), .rst(rst),
                    .ain1(aout49_8), .ain2(aout50_8), .ain3(aout51_8), .ain4(aout52_8),
                    .win1(wout48_9), .win2(wout48_10), .win3(wout48_11), .win4(wout48_12),
                    .aout1(aout49_12), .aout2(aout50_12), .aout3(aout51_12), .aout4(aout52_12),
                    .wout1(wout52_9), .wout2(wout52_10), .wout3(wout52_11), .wout4(wout52_12),
                    .sout11(sout49_9), .sout12(sout49_10), .sout13(sout49_11), .sout14(sout49_12),
                    .sout21(sout50_9), .sout22(sout50_10), .sout23(sout50_11), .sout24(sout50_12),
                    .sout31(sout51_9), .sout32(sout51_10), .sout33(sout51_11), .sout34(sout51_12),
                    .sout41(sout52_9), .sout42(sout52_10), .sout43(sout52_11), .sout44(sout52_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_13_4 (.clk(clk), .rst(rst),
                    .ain1(aout49_12), .ain2(aout50_12), .ain3(aout51_12), .ain4(aout52_12),
                    .win1(wout48_13), .win2(wout48_14), .win3(wout48_15), .win4(wout48_16),
                    .aout1(aout49_16), .aout2(aout50_16), .aout3(aout51_16), .aout4(aout52_16),
                    .wout1(wout52_13), .wout2(wout52_14), .wout3(wout52_15), .wout4(wout52_16),
                    .sout11(sout49_13), .sout12(sout49_14), .sout13(sout49_15), .sout14(sout49_16),
                    .sout21(sout50_13), .sout22(sout50_14), .sout23(sout50_15), .sout24(sout50_16),
                    .sout31(sout51_13), .sout32(sout51_14), .sout33(sout51_15), .sout34(sout51_16),
                    .sout41(sout52_13), .sout42(sout52_14), .sout43(sout52_15), .sout44(sout52_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_13_5 (.clk(clk), .rst(rst),
                    .ain1(aout49_16), .ain2(aout50_16), .ain3(aout51_16), .ain4(aout52_16),
                    .win1(wout48_17), .win2(wout48_18), .win3(wout48_19), .win4(wout48_20),
                    .aout1(aout49_20), .aout2(aout50_20), .aout3(aout51_20), .aout4(aout52_20),
                    .wout1(wout52_17), .wout2(wout52_18), .wout3(wout52_19), .wout4(wout52_20),
                    .sout11(sout49_17), .sout12(sout49_18), .sout13(sout49_19), .sout14(sout49_20),
                    .sout21(sout50_17), .sout22(sout50_18), .sout23(sout50_19), .sout24(sout50_20),
                    .sout31(sout51_17), .sout32(sout51_18), .sout33(sout51_19), .sout34(sout51_20),
                    .sout41(sout52_17), .sout42(sout52_18), .sout43(sout52_19), .sout44(sout52_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_13_6 (.clk(clk), .rst(rst),
                    .ain1(aout49_20), .ain2(aout50_20), .ain3(aout51_20), .ain4(aout52_20),
                    .win1(wout48_21), .win2(wout48_22), .win3(wout48_23), .win4(wout48_24),
                    .aout1(aout49_24), .aout2(aout50_24), .aout3(aout51_24), .aout4(aout52_24),
                    .wout1(wout52_21), .wout2(wout52_22), .wout3(wout52_23), .wout4(wout52_24),
                    .sout11(sout49_21), .sout12(sout49_22), .sout13(sout49_23), .sout14(sout49_24),
                    .sout21(sout50_21), .sout22(sout50_22), .sout23(sout50_23), .sout24(sout50_24),
                    .sout31(sout51_21), .sout32(sout51_22), .sout33(sout51_23), .sout34(sout51_24),
                    .sout41(sout52_21), .sout42(sout52_22), .sout43(sout52_23), .sout44(sout52_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_13_7 (.clk(clk), .rst(rst),
                    .ain1(aout49_24), .ain2(aout50_24), .ain3(aout51_24), .ain4(aout52_24),
                    .win1(wout48_25), .win2(wout48_26), .win3(wout48_27), .win4(wout48_28),
                    .aout1(aout49_28), .aout2(aout50_28), .aout3(aout51_28), .aout4(aout52_28),
                    .wout1(wout52_25), .wout2(wout52_26), .wout3(wout52_27), .wout4(wout52_28),
                    .sout11(sout49_25), .sout12(sout49_26), .sout13(sout49_27), .sout14(sout49_28),
                    .sout21(sout50_25), .sout22(sout50_26), .sout23(sout50_27), .sout24(sout50_28),
                    .sout31(sout51_25), .sout32(sout51_26), .sout33(sout51_27), .sout34(sout51_28),
                    .sout41(sout52_25), .sout42(sout52_26), .sout43(sout52_27), .sout44(sout52_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_13_8 (.clk(clk), .rst(rst),
                    .ain1(aout49_28), .ain2(aout50_28), .ain3(aout51_28), .ain4(aout52_28),
                    .win1(wout48_29), .win2(wout48_30), .win3(wout48_31), .win4(wout48_32),
                    .aout1(aout49_32), .aout2(aout50_32), .aout3(aout51_32), .aout4(aout52_32),
                    .wout1(wout52_29), .wout2(wout52_30), .wout3(wout52_31), .wout4(wout52_32),
                    .sout11(sout49_29), .sout12(sout49_30), .sout13(sout49_31), .sout14(sout49_32),
                    .sout21(sout50_29), .sout22(sout50_30), .sout23(sout50_31), .sout24(sout50_32),
                    .sout31(sout51_29), .sout32(sout51_30), .sout33(sout51_31), .sout34(sout51_32),
                    .sout41(sout52_29), .sout42(sout52_30), .sout43(sout52_31), .sout44(sout52_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_13_9 (.clk(clk), .rst(rst),
                    .ain1(aout49_32), .ain2(aout50_32), .ain3(aout51_32), .ain4(aout52_32),
                    .win1(wout48_33), .win2(wout48_34), .win3(wout48_35), .win4(wout48_36),
                    .aout1(aout49_36), .aout2(aout50_36), .aout3(aout51_36), .aout4(aout52_36),
                    .wout1(wout52_33), .wout2(wout52_34), .wout3(wout52_35), .wout4(wout52_36),
                    .sout11(sout49_33), .sout12(sout49_34), .sout13(sout49_35), .sout14(sout49_36),
                    .sout21(sout50_33), .sout22(sout50_34), .sout23(sout50_35), .sout24(sout50_36),
                    .sout31(sout51_33), .sout32(sout51_34), .sout33(sout51_35), .sout34(sout51_36),
                    .sout41(sout52_33), .sout42(sout52_34), .sout43(sout52_35), .sout44(sout52_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_13_10 (.clk(clk), .rst(rst),
                    .ain1(aout49_36), .ain2(aout50_36), .ain3(aout51_36), .ain4(aout52_36),
                    .win1(wout48_37), .win2(wout48_38), .win3(wout48_39), .win4(wout48_40),
                    .aout1(aout49_40), .aout2(aout50_40), .aout3(aout51_40), .aout4(aout52_40),
                    .wout1(wout52_37), .wout2(wout52_38), .wout3(wout52_39), .wout4(wout52_40),
                    .sout11(sout49_37), .sout12(sout49_38), .sout13(sout49_39), .sout14(sout49_40),
                    .sout21(sout50_37), .sout22(sout50_38), .sout23(sout50_39), .sout24(sout50_40),
                    .sout31(sout51_37), .sout32(sout51_38), .sout33(sout51_39), .sout34(sout51_40),
                    .sout41(sout52_37), .sout42(sout52_38), .sout43(sout52_39), .sout44(sout52_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_13_11 (.clk(clk), .rst(rst),
                    .ain1(aout49_40), .ain2(aout50_40), .ain3(aout51_40), .ain4(aout52_40),
                    .win1(wout48_41), .win2(wout48_42), .win3(wout48_43), .win4(wout48_44),
                    .aout1(aout49_44), .aout2(aout50_44), .aout3(aout51_44), .aout4(aout52_44),
                    .wout1(wout52_41), .wout2(wout52_42), .wout3(wout52_43), .wout4(wout52_44),
                    .sout11(sout49_41), .sout12(sout49_42), .sout13(sout49_43), .sout14(sout49_44),
                    .sout21(sout50_41), .sout22(sout50_42), .sout23(sout50_43), .sout24(sout50_44),
                    .sout31(sout51_41), .sout32(sout51_42), .sout33(sout51_43), .sout34(sout51_44),
                    .sout41(sout52_41), .sout42(sout52_42), .sout43(sout52_43), .sout44(sout52_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_13_12 (.clk(clk), .rst(rst),
                    .ain1(aout49_44), .ain2(aout50_44), .ain3(aout51_44), .ain4(aout52_44),
                    .win1(wout48_45), .win2(wout48_46), .win3(wout48_47), .win4(wout48_48),
                    .aout1(aout49_48), .aout2(aout50_48), .aout3(aout51_48), .aout4(aout52_48),
                    .wout1(wout52_45), .wout2(wout52_46), .wout3(wout52_47), .wout4(wout52_48),
                    .sout11(sout49_45), .sout12(sout49_46), .sout13(sout49_47), .sout14(sout49_48),
                    .sout21(sout50_45), .sout22(sout50_46), .sout23(sout50_47), .sout24(sout50_48),
                    .sout31(sout51_45), .sout32(sout51_46), .sout33(sout51_47), .sout34(sout51_48),
                    .sout41(sout52_45), .sout42(sout52_46), .sout43(sout52_47), .sout44(sout52_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_13_13 (.clk(clk), .rst(rst),
                    .ain1(aout49_48), .ain2(aout50_48), .ain3(aout51_48), .ain4(aout52_48),
                    .win1(wout48_49), .win2(wout48_50), .win3(wout48_51), .win4(wout48_52),
                    .aout1(aout49_52), .aout2(aout50_52), .aout3(aout51_52), .aout4(aout52_52),
                    .wout1(wout52_49), .wout2(wout52_50), .wout3(wout52_51), .wout4(wout52_52),
                    .sout11(sout49_49), .sout12(sout49_50), .sout13(sout49_51), .sout14(sout49_52),
                    .sout21(sout50_49), .sout22(sout50_50), .sout23(sout50_51), .sout24(sout50_52),
                    .sout31(sout51_49), .sout32(sout51_50), .sout33(sout51_51), .sout34(sout51_52),
                    .sout41(sout52_49), .sout42(sout52_50), .sout43(sout52_51), .sout44(sout52_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_13_14 (.clk(clk), .rst(rst),
                    .ain1(aout49_52), .ain2(aout50_52), .ain3(aout51_52), .ain4(aout52_52),
                    .win1(wout48_53), .win2(wout48_54), .win3(wout48_55), .win4(wout48_56),
                    .aout1(aout49_56), .aout2(aout50_56), .aout3(aout51_56), .aout4(aout52_56),
                    .wout1(wout52_53), .wout2(wout52_54), .wout3(wout52_55), .wout4(wout52_56),
                    .sout11(sout49_53), .sout12(sout49_54), .sout13(sout49_55), .sout14(sout49_56),
                    .sout21(sout50_53), .sout22(sout50_54), .sout23(sout50_55), .sout24(sout50_56),
                    .sout31(sout51_53), .sout32(sout51_54), .sout33(sout51_55), .sout34(sout51_56),
                    .sout41(sout52_53), .sout42(sout52_54), .sout43(sout52_55), .sout44(sout52_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_13_15 (.clk(clk), .rst(rst),
                    .ain1(aout49_56), .ain2(aout50_56), .ain3(aout51_56), .ain4(aout52_56),
                    .win1(wout48_57), .win2(wout48_58), .win3(wout48_59), .win4(wout48_60),
                    .aout1(aout49_60), .aout2(aout50_60), .aout3(aout51_60), .aout4(aout52_60),
                    .wout1(wout52_57), .wout2(wout52_58), .wout3(wout52_59), .wout4(wout52_60),
                    .sout11(sout49_57), .sout12(sout49_58), .sout13(sout49_59), .sout14(sout49_60),
                    .sout21(sout50_57), .sout22(sout50_58), .sout23(sout50_59), .sout24(sout50_60),
                    .sout31(sout51_57), .sout32(sout51_58), .sout33(sout51_59), .sout34(sout51_60),
                    .sout41(sout52_57), .sout42(sout52_58), .sout43(sout52_59), .sout44(sout52_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_13_16 (.clk(clk), .rst(rst),
                    .ain1(aout49_60), .ain2(aout50_60), .ain3(aout51_60), .ain4(aout52_60),
                    .win1(wout48_61), .win2(wout48_62), .win3(wout48_63), .win4(wout48_64),
                    .aout1(aout49_64), .aout2(aout50_64), .aout3(aout51_64), .aout4(aout52_64),
                    .wout1(wout52_61), .wout2(wout52_62), .wout3(wout52_63), .wout4(wout52_64),
                    .sout11(sout49_61), .sout12(sout49_62), .sout13(sout49_63), .sout14(sout49_64),
                    .sout21(sout50_61), .sout22(sout50_62), .sout23(sout50_63), .sout24(sout50_64),
                    .sout31(sout51_61), .sout32(sout51_62), .sout33(sout51_63), .sout34(sout51_64),
                    .sout41(sout52_61), .sout42(sout52_62), .sout43(sout52_63), .sout44(sout52_64)
                    ); //4x4 MAC array
    
    
    //row14
    mac_array_4x4 mac_array_4x4_14_1 (.clk(clk), .rst(rst),
                    .ain1(ain53), .ain2(ain54), .ain3(ain55), .ain4(ain56),
                    .win1(wout52_1), .win2(wout52_2), .win3(wout52_3), .win4(wout52_4),
                    .aout1(aout53_4), .aout2(aout54_4), .aout3(aout55_4), .aout4(aout56_4),
                    .wout1(wout56_1), .wout2(wout56_2), .wout3(wout56_3), .wout4(wout56_4),
                    .sout11(sout53_1), .sout12(sout53_2), .sout13(sout53_3), .sout14(sout53_4),
                    .sout21(sout54_1), .sout22(sout54_2), .sout23(sout54_3), .sout24(sout54_4),
                    .sout31(sout55_1), .sout32(sout55_2), .sout33(sout55_3), .sout34(sout55_4),
                    .sout41(sout56_1), .sout42(sout56_2), .sout43(sout56_3), .sout44(sout56_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_14_2 (.clk(clk), .rst(rst),
                    .ain1(aout53_4), .ain2(aout54_4), .ain3(aout55_4), .ain4(aout56_4),
                    .win1(wout52_5), .win2(wout52_6), .win3(wout52_7), .win4(wout52_8),
                    .aout1(aout53_8), .aout2(aout54_8), .aout3(aout55_8), .aout4(aout56_8),
                    .wout1(wout56_5), .wout2(wout56_6), .wout3(wout56_7), .wout4(wout56_8),
                    .sout11(sout53_5), .sout12(sout53_6), .sout13(sout53_7), .sout14(sout53_8),
                    .sout21(sout54_5), .sout22(sout54_6), .sout23(sout54_7), .sout24(sout54_8),
                    .sout31(sout55_5), .sout32(sout55_6), .sout33(sout55_7), .sout34(sout55_8),
                    .sout41(sout56_5), .sout42(sout56_6), .sout43(sout56_7), .sout44(sout56_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_14_3 (.clk(clk), .rst(rst),
                    .ain1(aout53_8), .ain2(aout54_8), .ain3(aout55_8), .ain4(aout56_8),
                    .win1(wout52_9), .win2(wout52_10), .win3(wout52_11), .win4(wout52_12),
                    .aout1(aout53_12), .aout2(aout54_12), .aout3(aout55_12), .aout4(aout56_12),
                    .wout1(wout56_9), .wout2(wout56_10), .wout3(wout56_11), .wout4(wout56_12),
                    .sout11(sout53_9), .sout12(sout53_10), .sout13(sout53_11), .sout14(sout53_12),
                    .sout21(sout54_9), .sout22(sout54_10), .sout23(sout54_11), .sout24(sout54_12),
                    .sout31(sout55_9), .sout32(sout55_10), .sout33(sout55_11), .sout34(sout55_12),
                    .sout41(sout56_9), .sout42(sout56_10), .sout43(sout56_11), .sout44(sout56_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14_4 (.clk(clk), .rst(rst),
                    .ain1(aout53_12), .ain2(aout54_12), .ain3(aout55_12), .ain4(aout56_12),
                    .win1(wout52_13), .win2(wout52_14), .win3(wout52_15), .win4(wout52_16),
                    .aout1(aout53_16), .aout2(aout54_16), .aout3(aout55_16), .aout4(aout56_16),
                    .wout1(wout56_13), .wout2(wout56_14), .wout3(wout56_15), .wout4(wout56_16),
                    .sout11(sout53_13), .sout12(sout53_14), .sout13(sout53_15), .sout14(sout53_16),
                    .sout21(sout54_13), .sout22(sout54_14), .sout23(sout54_15), .sout24(sout54_16),
                    .sout31(sout55_13), .sout32(sout55_14), .sout33(sout55_15), .sout34(sout55_16),
                    .sout41(sout56_13), .sout42(sout56_14), .sout43(sout56_15), .sout44(sout56_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14_5 (.clk(clk), .rst(rst),
                    .ain1(aout53_16), .ain2(aout54_16), .ain3(aout55_16), .ain4(aout56_16),
                    .win1(wout52_17), .win2(wout52_18), .win3(wout52_19), .win4(wout52_20),
                    .aout1(aout53_20), .aout2(aout54_20), .aout3(aout55_20), .aout4(aout56_20),
                    .wout1(wout56_17), .wout2(wout56_18), .wout3(wout56_19), .wout4(wout56_20),
                    .sout11(sout53_17), .sout12(sout53_18), .sout13(sout53_19), .sout14(sout53_20),
                    .sout21(sout54_17), .sout22(sout54_18), .sout23(sout54_19), .sout24(sout54_20),
                    .sout31(sout55_17), .sout32(sout55_18), .sout33(sout55_19), .sout34(sout55_20),
                    .sout41(sout56_17), .sout42(sout56_18), .sout43(sout56_19), .sout44(sout56_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_14_6 (.clk(clk), .rst(rst),
                    .ain1(aout53_20), .ain2(aout54_20), .ain3(aout55_20), .ain4(aout56_20),
                    .win1(wout52_21), .win2(wout52_22), .win3(wout52_23), .win4(wout52_24),
                    .aout1(aout53_24), .aout2(aout54_24), .aout3(aout55_24), .aout4(aout56_24),
                    .wout1(wout56_21), .wout2(wout56_22), .wout3(wout56_23), .wout4(wout56_24),
                    .sout11(sout53_21), .sout12(sout53_22), .sout13(sout53_23), .sout14(sout53_24),
                    .sout21(sout54_21), .sout22(sout54_22), .sout23(sout54_23), .sout24(sout54_24),
                    .sout31(sout55_21), .sout32(sout55_22), .sout33(sout55_23), .sout34(sout55_24),
                    .sout41(sout56_21), .sout42(sout56_22), .sout43(sout56_23), .sout44(sout56_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14_7 (.clk(clk), .rst(rst),
                    .ain1(aout53_24), .ain2(aout54_24), .ain3(aout55_24), .ain4(aout56_24),
                    .win1(wout52_25), .win2(wout52_26), .win3(wout52_27), .win4(wout52_28),
                    .aout1(aout53_28), .aout2(aout54_28), .aout3(aout55_28), .aout4(aout56_28),
                    .wout1(wout56_25), .wout2(wout56_26), .wout3(wout56_27), .wout4(wout56_28),
                    .sout11(sout53_25), .sout12(sout53_26), .sout13(sout53_27), .sout14(sout53_28),
                    .sout21(sout54_25), .sout22(sout54_26), .sout23(sout54_27), .sout24(sout54_28),
                    .sout31(sout55_25), .sout32(sout55_26), .sout33(sout55_27), .sout34(sout55_28),
                    .sout41(sout56_25), .sout42(sout56_26), .sout43(sout56_27), .sout44(sout56_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_14_8 (.clk(clk), .rst(rst),
                    .ain1(aout53_28), .ain2(aout54_28), .ain3(aout55_28), .ain4(aout56_28),
                    .win1(wout52_29), .win2(wout52_30), .win3(wout52_31), .win4(wout52_32),
                    .aout1(aout53_32), .aout2(aout54_32), .aout3(aout55_32), .aout4(aout56_32),
                    .wout1(wout56_29), .wout2(wout56_30), .wout3(wout56_31), .wout4(wout56_32),
                    .sout11(sout53_29), .sout12(sout53_30), .sout13(sout53_31), .sout14(sout53_32),
                    .sout21(sout54_29), .sout22(sout54_30), .sout23(sout54_31), .sout24(sout54_32),
                    .sout31(sout55_29), .sout32(sout55_30), .sout33(sout55_31), .sout34(sout55_32),
                    .sout41(sout56_29), .sout42(sout56_30), .sout43(sout56_31), .sout44(sout56_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14_9 (.clk(clk), .rst(rst),
                    .ain1(aout53_32), .ain2(aout54_32), .ain3(aout55_32), .ain4(aout56_32),
                    .win1(wout52_33), .win2(wout52_34), .win3(wout52_35), .win4(wout52_36),
                    .aout1(aout53_36), .aout2(aout54_36), .aout3(aout55_36), .aout4(aout56_36),
                    .wout1(wout56_33), .wout2(wout56_34), .wout3(wout56_35), .wout4(wout56_36),
                    .sout11(sout53_33), .sout12(sout53_34), .sout13(sout53_35), .sout14(sout53_36),
                    .sout21(sout54_33), .sout22(sout54_34), .sout23(sout54_35), .sout24(sout54_36),
                    .sout31(sout55_33), .sout32(sout55_34), .sout33(sout55_35), .sout34(sout55_36),
                    .sout41(sout56_33), .sout42(sout56_34), .sout43(sout56_35), .sout44(sout56_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14_10 (.clk(clk), .rst(rst),
                    .ain1(aout53_36), .ain2(aout54_36), .ain3(aout55_36), .ain4(aout56_36),
                    .win1(wout52_37), .win2(wout52_38), .win3(wout52_39), .win4(wout52_40),
                    .aout1(aout53_40), .aout2(aout54_40), .aout3(aout55_40), .aout4(aout56_40),
                    .wout1(wout56_37), .wout2(wout56_38), .wout3(wout56_39), .wout4(wout56_40),
                    .sout11(sout53_37), .sout12(sout53_38), .sout13(sout53_39), .sout14(sout53_40),
                    .sout21(sout54_37), .sout22(sout54_38), .sout23(sout54_39), .sout24(sout54_40),
                    .sout31(sout55_37), .sout32(sout55_38), .sout33(sout55_39), .sout34(sout55_40),
                    .sout41(sout56_37), .sout42(sout56_38), .sout43(sout56_39), .sout44(sout56_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14_11 (.clk(clk), .rst(rst),
                    .ain1(aout53_40), .ain2(aout54_40), .ain3(aout55_40), .ain4(aout56_40),
                    .win1(wout52_41), .win2(wout52_42), .win3(wout52_43), .win4(wout52_44),
                    .aout1(aout53_44), .aout2(aout54_44), .aout3(aout55_44), .aout4(aout56_44),
                    .wout1(wout56_41), .wout2(wout56_42), .wout3(wout56_43), .wout4(wout56_44),
                    .sout11(sout53_41), .sout12(sout53_42), .sout13(sout53_43), .sout14(sout53_44),
                    .sout21(sout54_41), .sout22(sout54_42), .sout23(sout54_43), .sout24(sout54_44),
                    .sout31(sout55_41), .sout32(sout55_42), .sout33(sout55_43), .sout34(sout55_44),
                    .sout41(sout56_41), .sout42(sout56_42), .sout43(sout56_43), .sout44(sout56_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14_12 (.clk(clk), .rst(rst),
                    .ain1(aout53_44), .ain2(aout54_44), .ain3(aout55_44), .ain4(aout56_44),
                    .win1(wout52_45), .win2(wout52_46), .win3(wout52_47), .win4(wout52_48),
                    .aout1(aout53_48), .aout2(aout54_48), .aout3(aout55_48), .aout4(aout56_48),
                    .wout1(wout56_45), .wout2(wout56_46), .wout3(wout56_47), .wout4(wout56_48),
                    .sout11(sout53_45), .sout12(sout53_46), .sout13(sout53_47), .sout14(sout53_48),
                    .sout21(sout54_45), .sout22(sout54_46), .sout23(sout54_47), .sout24(sout54_48),
                    .sout31(sout55_45), .sout32(sout55_46), .sout33(sout55_47), .sout34(sout55_48),
                    .sout41(sout56_45), .sout42(sout56_46), .sout43(sout56_47), .sout44(sout56_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14_13 (.clk(clk), .rst(rst),
                    .ain1(aout53_48), .ain2(aout54_48), .ain3(aout55_48), .ain4(aout56_48),
                    .win1(wout52_49), .win2(wout52_50), .win3(wout52_51), .win4(wout52_52),
                    .aout1(aout53_52), .aout2(aout54_52), .aout3(aout55_52), .aout4(aout56_52),
                    .wout1(wout56_49), .wout2(wout56_50), .wout3(wout56_51), .wout4(wout56_52),
                    .sout11(sout53_49), .sout12(sout53_50), .sout13(sout53_51), .sout14(sout53_52),
                    .sout21(sout54_49), .sout22(sout54_50), .sout23(sout54_51), .sout24(sout54_52),
                    .sout31(sout55_49), .sout32(sout55_50), .sout33(sout55_51), .sout34(sout55_52),
                    .sout41(sout56_49), .sout42(sout56_50), .sout43(sout56_51), .sout44(sout56_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14_14 (.clk(clk), .rst(rst),
                    .ain1(aout53_52), .ain2(aout54_52), .ain3(aout55_52), .ain4(aout56_52),
                    .win1(wout52_53), .win2(wout52_54), .win3(wout52_55), .win4(wout52_56),
                    .aout1(aout53_56), .aout2(aout54_56), .aout3(aout55_56), .aout4(aout56_56),
                    .wout1(wout56_53), .wout2(wout56_54), .wout3(wout56_55), .wout4(wout56_56),
                    .sout11(sout53_53), .sout12(sout53_54), .sout13(sout53_55), .sout14(sout53_56),
                    .sout21(sout54_53), .sout22(sout54_54), .sout23(sout54_55), .sout24(sout54_56),
                    .sout31(sout55_53), .sout32(sout55_54), .sout33(sout55_55), .sout34(sout55_56),
                    .sout41(sout56_53), .sout42(sout56_54), .sout43(sout56_55), .sout44(sout56_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_14_15 (.clk(clk), .rst(rst),
                    .ain1(aout53_56), .ain2(aout54_56), .ain3(aout55_56), .ain4(aout56_56),
                    .win1(wout52_57), .win2(wout52_58), .win3(wout52_59), .win4(wout52_60),
                    .aout1(aout53_60), .aout2(aout54_60), .aout3(aout55_60), .aout4(aout56_60),
                    .wout1(wout52_57), .wout2(wout52_58), .wout3(wout52_59), .wout4(wout52_60),
                    .sout11(sout53_57), .sout12(sout53_58), .sout13(sout53_59), .sout14(sout53_60),
                    .sout21(sout54_57), .sout22(sout54_58), .sout23(sout54_59), .sout24(sout54_60),
                    .sout31(sout55_57), .sout32(sout55_58), .sout33(sout55_59), .sout34(sout55_60),
                    .sout41(sout56_57), .sout42(sout56_58), .sout43(sout56_59), .sout44(sout56_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_14_16 (.clk(clk), .rst(rst),
                    .ain1(aout53_60), .ain2(aout54_60), .ain3(aout55_60), .ain4(aout56_60),
                    .win1(wout52_61), .win2(wout52_62), .win3(wout52_63), .win4(wout52_64),
                    .aout1(aout53_64), .aout2(aout54_64), .aout3(aout55_64), .aout4(aout56_64),
                    .wout1(wout56_61), .wout2(wout56_62), .wout3(wout56_63), .wout4(wout56_64),
                    .sout11(sout53_61), .sout12(sout53_62), .sout13(sout53_63), .sout14(sout53_64),
                    .sout21(sout54_61), .sout22(sout54_62), .sout23(sout54_63), .sout24(sout54_64),
                    .sout31(sout55_61), .sout32(sout55_62), .sout33(sout55_63), .sout34(sout55_64),
                    .sout41(sout56_61), .sout42(sout56_62), .sout43(sout56_63), .sout44(sout56_64)
                    ); //4x4 MAC array
                    
                    
    //row15
    mac_array_4x4 mac_array_4x4_15_1 (.clk(clk), .rst(rst),
                    .ain1(ain57), .ain2(ain58), .ain3(ain59), .ain4(ain60),
                    .win1(wout56_1), .win2(wout56_2), .win3(wout56_3), .win4(wout56_4),
                    .aout1(aout57_4), .aout2(aout58_4), .aout3(aout59_4), .aout4(aout60_4),
                    .wout1(wout60_1), .wout2(wout60_2), .wout3(wout60_3), .wout4(wout60_4),
                    .sout11(sout57_1), .sout12(sout57_2), .sout13(sout57_3), .sout14(sout57_4),
                    .sout21(sout58_1), .sout22(sout58_2), .sout23(sout58_3), .sout24(sout58_4),
                    .sout31(sout59_1), .sout32(sout59_2), .sout33(sout59_3), .sout34(sout59_4),
                    .sout41(sout60_1), .sout42(sout60_2), .sout43(sout60_3), .sout44(sout60_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_15_2 (.clk(clk), .rst(rst),
                    .ain1(aout57_4), .ain2(aout58_4), .ain3(aout59_4), .ain4(aout60_4),
                    .win1(wout56_5), .win2(wout56_6), .win3(wout56_7), .win4(wout56_8),
                    .aout1(aout57_8), .aout2(aout58_8), .aout3(aout59_8), .aout4(aout60_8),
                    .wout1(wout60_5), .wout2(wout60_6), .wout3(wout60_7), .wout4(wout60_8),
                    .sout11(sout57_5), .sout12(sout57_6), .sout13(sout57_7), .sout14(sout57_8),
                    .sout21(sout58_5), .sout22(sout58_6), .sout23(sout58_7), .sout24(sout58_8),
                    .sout31(sout59_5), .sout32(sout59_6), .sout33(sout59_7), .sout34(sout59_8),
                    .sout41(sout60_5), .sout42(sout60_6), .sout43(sout60_7), .sout44(sout60_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_15_3 (.clk(clk), .rst(rst),
                    .ain1(aout57_8), .ain2(aout58_8), .ain3(aout59_8), .ain4(aout60_8),
                    .win1(wout56_9), .win2(wout56_10), .win3(wout56_11), .win4(wout56_12),
                    .aout1(aout57_12), .aout2(aout58_12), .aout3(aout59_12), .aout4(aout60_12),
                    .wout1(wout60_9), .wout2(wout60_10), .wout3(wout60_11), .wout4(wout60_12),
                    .sout11(sout57_9), .sout12(sout57_10), .sout13(sout57_11), .sout14(sout57_12),
                    .sout21(sout58_9), .sout22(sout58_10), .sout23(sout58_11), .sout24(sout58_12),
                    .sout31(sout59_9), .sout32(sout59_10), .sout33(sout59_11), .sout34(sout59_12),
                    .sout41(sout60_9), .sout42(sout60_10), .sout43(sout60_11), .sout44(sout60_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15_4 (.clk(clk), .rst(rst),
                    .ain1(aout57_12), .ain2(aout58_12), .ain3(aout59_12), .ain4(aout60_12),
                    .win1(wout56_13), .win2(wout56_14), .win3(wout56_15), .win4(wout56_16),
                    .aout1(aout57_16), .aout2(aout58_16), .aout3(aout59_16), .aout4(aout60_16),
                    .wout1(wout60_13), .wout2(wout60_14), .wout3(wout60_15), .wout4(wout60_16),
                    .sout11(sout57_13), .sout12(sout57_14), .sout13(sout57_15), .sout14(sout57_16),
                    .sout21(sout58_13), .sout22(sout58_14), .sout23(sout58_15), .sout24(sout58_16),
                    .sout31(sout59_13), .sout32(sout59_14), .sout33(sout59_15), .sout34(sout59_16),
                    .sout41(sout60_13), .sout42(sout60_14), .sout43(sout60_15), .sout44(sout60_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15_5 (.clk(clk), .rst(rst),
                    .ain1(aout57_16), .ain2(aout58_16), .ain3(aout59_16), .ain4(aout60_16),
                    .win1(wout56_17), .win2(wout56_18), .win3(wout56_19), .win4(wout56_20),
                    .aout1(aout57_20), .aout2(aout58_20), .aout3(aout59_20), .aout4(aout60_20),
                    .wout1(wout60_17), .wout2(wout60_18), .wout3(wout60_19), .wout4(wout60_20),
                    .sout11(sout57_17), .sout12(sout57_18), .sout13(sout57_19), .sout14(sout57_20),
                    .sout21(sout58_17), .sout22(sout58_18), .sout23(sout58_19), .sout24(sout58_20),
                    .sout31(sout59_17), .sout32(sout59_18), .sout33(sout59_19), .sout34(sout59_20),
                    .sout41(sout60_17), .sout42(sout60_18), .sout43(sout60_19), .sout44(sout60_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_15_6 (.clk(clk), .rst(rst),
                    .ain1(aout57_20), .ain2(aout58_20), .ain3(aout59_20), .ain4(aout60_20),
                    .win1(wout56_21), .win2(wout56_22), .win3(wout56_23), .win4(wout56_24),
                    .aout1(aout57_24), .aout2(aout58_24), .aout3(aout59_24), .aout4(aout60_24),
                    .wout1(wout60_21), .wout2(wout60_22), .wout3(wout60_23), .wout4(wout60_24),
                    .sout11(sout57_21), .sout12(sout57_22), .sout13(sout57_23), .sout14(sout57_24),
                    .sout21(sout58_21), .sout22(sout58_22), .sout23(sout58_23), .sout24(sout58_24),
                    .sout31(sout59_21), .sout32(sout59_22), .sout33(sout59_23), .sout34(sout59_24),
                    .sout41(sout60_21), .sout42(sout60_22), .sout43(sout60_23), .sout44(sout60_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15_7 (.clk(clk), .rst(rst),
                    .ain1(aout57_24), .ain2(aout58_24), .ain3(aout59_24), .ain4(aout60_24),
                    .win1(wout56_25), .win2(wout56_26), .win3(wout56_27), .win4(wout56_28),
                    .aout1(aout57_28), .aout2(aout58_28), .aout3(aout59_28), .aout4(aout60_28),
                    .wout1(wout60_25), .wout2(wout60_26), .wout3(wout60_27), .wout4(wout60_28),
                    .sout11(sout57_25), .sout12(sout57_26), .sout13(sout57_27), .sout14(sout57_28),
                    .sout21(sout58_25), .sout22(sout58_26), .sout23(sout58_27), .sout24(sout58_28),
                    .sout31(sout59_25), .sout32(sout59_26), .sout33(sout59_27), .sout34(sout59_28),
                    .sout41(sout60_25), .sout42(sout60_26), .sout43(sout60_27), .sout44(sout60_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_15_8 (.clk(clk), .rst(rst),
                    .ain1(aout57_28), .ain2(aout58_28), .ain3(aout59_28), .ain4(aout60_28),
                    .win1(wout56_29), .win2(wout56_30), .win3(wout56_31), .win4(wout56_32),
                    .aout1(aout57_32), .aout2(aout58_32), .aout3(aout59_32), .aout4(aout60_32),
                    .wout1(wout60_29), .wout2(wout60_30), .wout3(wout60_31), .wout4(wout60_32),
                    .sout11(sout57_29), .sout12(sout57_30), .sout13(sout57_31), .sout14(sout57_32),
                    .sout21(sout58_29), .sout22(sout58_30), .sout23(sout58_31), .sout24(sout58_32),
                    .sout31(sout59_29), .sout32(sout59_30), .sout33(sout59_31), .sout34(sout59_32),
                    .sout41(sout60_29), .sout42(sout60_30), .sout43(sout60_31), .sout44(sout60_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15_9 (.clk(clk), .rst(rst),
                    .ain1(aout57_32), .ain2(aout58_32), .ain3(aout59_32), .ain4(aout60_32),
                    .win1(wout56_33), .win2(wout56_34), .win3(wout56_35), .win4(wout56_36),
                    .aout1(aout57_36), .aout2(aout58_36), .aout3(aout59_36), .aout4(aout60_36),
                    .wout1(wout60_33), .wout2(wout60_34), .wout3(wout60_35), .wout4(wout60_36),
                    .sout11(sout57_33), .sout12(sout57_34), .sout13(sout57_35), .sout14(sout57_36),
                    .sout21(sout58_33), .sout22(sout58_34), .sout23(sout58_35), .sout24(sout58_36),
                    .sout31(sout59_33), .sout32(sout59_34), .sout33(sout59_35), .sout34(sout59_36),
                    .sout41(sout60_33), .sout42(sout60_34), .sout43(sout60_35), .sout44(sout60_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15_10 (.clk(clk), .rst(rst),
                    .ain1(aout57_36), .ain2(aout58_36), .ain3(aout59_36), .ain4(aout60_36),
                    .win1(wout56_37), .win2(wout56_38), .win3(wout56_39), .win4(wout56_40),
                    .aout1(aout57_40), .aout2(aout58_40), .aout3(aout59_40), .aout4(aout60_40),
                    .wout1(wout60_37), .wout2(wout60_38), .wout3(wout60_39), .wout4(wout60_40),
                    .sout11(sout57_37), .sout12(sout57_38), .sout13(sout57_39), .sout14(sout57_40),
                    .sout21(sout58_37), .sout22(sout58_38), .sout23(sout58_39), .sout24(sout58_40),
                    .sout31(sout59_37), .sout32(sout59_38), .sout33(sout59_39), .sout34(sout59_40),
                    .sout41(sout60_37), .sout42(sout60_38), .sout43(sout60_39), .sout44(sout60_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15_11 (.clk(clk), .rst(rst),
                    .ain1(aout57_40), .ain2(aout58_40), .ain3(aout59_40), .ain4(aout60_40),
                    .win1(wout56_41), .win2(wout56_42), .win3(wout56_43), .win4(wout56_44),
                    .aout1(aout57_44), .aout2(aout58_44), .aout3(aout59_44), .aout4(aout60_44),
                    .wout1(wout60_41), .wout2(wout60_42), .wout3(wout60_43), .wout4(wout60_44),
                    .sout11(sout57_41), .sout12(sout57_42), .sout13(sout57_43), .sout14(sout57_44),
                    .sout21(sout58_41), .sout22(sout58_42), .sout23(sout58_43), .sout24(sout58_44),
                    .sout31(sout59_41), .sout32(sout59_42), .sout33(sout59_43), .sout34(sout59_44),
                    .sout41(sout60_41), .sout42(sout60_42), .sout43(sout60_43), .sout44(sout60_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15_12 (.clk(clk), .rst(rst),
                    .ain1(aout57_44), .ain2(aout58_44), .ain3(aout59_44), .ain4(aout60_44),
                    .win1(wout56_45), .win2(wout56_46), .win3(wout56_47), .win4(wout56_48),
                    .aout1(aout57_48), .aout2(aout58_48), .aout3(aout59_48), .aout4(aout60_48),
                    .wout1(wout60_45), .wout2(wout60_46), .wout3(wout60_47), .wout4(wout60_48),
                    .sout11(sout57_45), .sout12(sout57_46), .sout13(sout57_47), .sout14(sout57_48),
                    .sout21(sout58_45), .sout22(sout58_46), .sout23(sout58_47), .sout24(sout58_48),
                    .sout31(sout59_45), .sout32(sout59_46), .sout33(sout59_47), .sout34(sout59_48),
                    .sout41(sout60_45), .sout42(sout60_46), .sout43(sout60_47), .sout44(sout60_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15_13 (.clk(clk), .rst(rst),
                    .ain1(aout57_48), .ain2(aout58_48), .ain3(aout59_48), .ain4(aout60_48),
                    .win1(wout56_49), .win2(wout56_50), .win3(wout56_51), .win4(wout56_52),
                    .aout1(aout57_52), .aout2(aout58_52), .aout3(aout59_52), .aout4(aout60_52),
                    .wout1(wout60_49), .wout2(wout60_50), .wout3(wout60_51), .wout4(wout60_52),
                    .sout11(sout57_49), .sout12(sout57_50), .sout13(sout57_51), .sout14(sout57_52),
                    .sout21(sout58_49), .sout22(sout58_50), .sout23(sout58_51), .sout24(sout58_52),
                    .sout31(sout59_49), .sout32(sout59_50), .sout33(sout59_51), .sout34(sout59_52),
                    .sout41(sout60_49), .sout42(sout60_50), .sout43(sout60_51), .sout44(sout60_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15_14 (.clk(clk), .rst(rst),
                    .ain1(aout57_52), .ain2(aout58_52), .ain3(aout59_52), .ain4(aout60_52),
                    .win1(wout56_53), .win2(wout56_54), .win3(wout56_55), .win4(wout56_56),
                    .aout1(aout57_56), .aout2(aout58_56), .aout3(aout59_56), .aout4(aout60_56),
                    .wout1(wout60_53), .wout2(wout60_54), .wout3(wout60_55), .wout4(wout60_56),
                    .sout11(sout57_53), .sout12(sout57_54), .sout13(sout57_55), .sout14(sout57_56),
                    .sout21(sout58_53), .sout22(sout58_54), .sout23(sout58_55), .sout24(sout58_56),
                    .sout31(sout59_53), .sout32(sout59_54), .sout33(sout59_55), .sout34(sout59_56),
                    .sout41(sout60_53), .sout42(sout60_54), .sout43(sout60_55), .sout44(sout60_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_15_15 (.clk(clk), .rst(rst),
                    .ain1(aout57_56), .ain2(aout58_56), .ain3(aout59_56), .ain4(aout60_56),
                    .win1(wout56_57), .win2(wout56_58), .win3(wout56_59), .win4(wout56_60),
                    .aout1(aout57_60), .aout2(aout58_60), .aout3(aout59_60), .aout4(aout60_60),
                    .wout1(wout60_57), .wout2(wout60_58), .wout3(wout60_59), .wout4(wout60_60),
                    .sout11(sout57_57), .sout12(sout57_58), .sout13(sout57_59), .sout14(sout57_60),
                    .sout21(sout58_57), .sout22(sout58_58), .sout23(sout58_59), .sout24(sout58_60),
                    .sout31(sout59_57), .sout32(sout59_58), .sout33(sout59_59), .sout34(sout59_60),
                    .sout41(sout60_57), .sout42(sout60_58), .sout43(sout60_59), .sout44(sout60_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_15_16 (.clk(clk), .rst(rst),
                    .ain1(aout57_60), .ain2(aout58_60), .ain3(aout59_60), .ain4(aout60_60),
                    .win1(wout56_61), .win2(wout56_62), .win3(wout56_63), .win4(wout56_64),
                    .aout1(aout57_64), .aout2(aout58_64), .aout3(aout59_64), .aout4(aout60_64),
                    .wout1(wout60_61), .wout2(wout60_62), .wout3(wout60_63), .wout4(wout60_64),
                    .sout11(sout57_61), .sout12(sout57_62), .sout13(sout57_63), .sout14(sout57_64),
                    .sout21(sout58_61), .sout22(sout58_62), .sout23(sout58_63), .sout24(sout58_64),
                    .sout31(sout59_61), .sout32(sout59_62), .sout33(sout59_63), .sout34(sout59_64),
                    .sout41(sout60_61), .sout42(sout60_62), .sout43(sout60_63), .sout44(sout60_64)
                    ); //4x4 MAC array
                    
               
    //row16
    mac_array_4x4 mac_array_4x4_16_1 (.clk(clk), .rst(rst),
                    .ain1(ain61), .ain2(ain62), .ain3(ain63), .ain4(ain64),
                    .win1(wout60_1), .win2(wout60_2), .win3(wout60_3), .win4(wout60_4),
                    .aout1(aout61_4), .aout2(aout62_4), .aout3(aout63_4), .aout4(aout64_4),
                    .wout1(wout60_1), .wout2(wout60_2), .wout3(wout60_3), .wout4(wout60_4),
                    .sout11(sout57_1), .sout12(sout57_2), .sout13(sout57_3), .sout14(sout57_4),
                    .sout21(sout58_1), .sout22(sout58_2), .sout23(sout58_3), .sout24(sout58_4),
                    .sout31(sout59_1), .sout32(sout59_2), .sout33(sout59_3), .sout34(sout59_4),
                    .sout41(sout60_1), .sout42(sout60_2), .sout43(sout60_3), .sout44(sout60_4)
                    ); //4x4 MAC array
                    
  
    mac_array_4x4 mac_array_4x4_16_2 (.clk(clk), .rst(rst),
                    .ain1(aout61_4), .ain2(aout62_4), .ain3(aout63_4), .ain4(aout64_4),
                    .win1(wout60_5), .win2(wout60_6), .win3(wout60_7), .win4(wout60_8),
                    .aout1(aout61_8), .aout2(aout62_8), .aout3(aout63_8), .aout4(aout64_8),
                    .wout1(wout64_5), .wout2(wout64_6), .wout3(wout64_7), .wout4(wout64_8),
                    .sout11(sout61_5), .sout12(sout61_6), .sout13(sout61_7), .sout14(sout61_8),
                    .sout21(sout62_5), .sout22(sout62_6), .sout23(sout62_7), .sout24(sout62_8),
                    .sout31(sout63_5), .sout32(sout63_6), .sout33(sout63_7), .sout34(sout63_8),
                    .sout41(sout64_5), .sout42(sout64_6), .sout43(sout64_7), .sout44(sout64_8)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_16_3 (.clk(clk), .rst(rst),
                    .ain1(aout61_8), .ain2(aout62_8), .ain3(aout63_8), .ain4(aout64_8),
                    .win1(wout60_9), .win2(wout60_10), .win3(wout60_11), .win4(wout60_12),
                    .aout1(aout61_12), .aout2(aout62_12), .aout3(aout63_12), .aout4(aout64_12),
                    .wout1(wout64_9), .wout2(wout64_10), .wout3(wout64_11), .wout4(wout64_12),
                    .sout11(sout61_9), .sout12(sout61_10), .sout13(sout61_11), .sout14(sout61_12),
                    .sout21(sout62_9), .sout22(sout62_10), .sout23(sout62_11), .sout24(sout62_12),
                    .sout31(sout63_9), .sout32(sout63_10), .sout33(sout63_11), .sout34(sout63_12),
                    .sout41(sout64_9), .sout42(sout64_10), .sout43(sout64_11), .sout44(sout64_12)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16_4 (.clk(clk), .rst(rst),
                    .ain1(aout61_12), .ain2(aout62_12), .ain3(aout63_12), .ain4(aout64_12),
                    .win1(wout60_13), .win2(wout60_14), .win3(wout60_15), .win4(wout60_16),
                    .aout1(aout61_16), .aout2(aout62_16), .aout3(aout63_16), .aout4(aout64_16),
                    .wout1(wout64_13), .wout2(wout64_14), .wout3(wout64_15), .wout4(wout64_16),
                    .sout11(sout61_13), .sout12(sout61_14), .sout13(sout61_15), .sout14(sout61_16),
                    .sout21(sout62_13), .sout22(sout62_14), .sout23(sout62_15), .sout24(sout62_16),
                    .sout31(sout63_13), .sout32(sout63_14), .sout33(sout63_15), .sout34(sout63_16),
                    .sout41(sout64_13), .sout42(sout64_14), .sout43(sout64_15), .sout44(sout64_16)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16_5 (.clk(clk), .rst(rst),
                    .ain1(aout61_16), .ain2(aout62_16), .ain3(aout63_16), .ain4(aout64_16),
                    .win1(wout60_17), .win2(wout60_18), .win3(wout60_19), .win4(wout60_20),
                    .aout1(aout61_20), .aout2(aout62_20), .aout3(aout63_20), .aout4(aout64_20),
                    .wout1(wout64_17), .wout2(wout64_18), .wout3(wout64_19), .wout4(wout64_20),
                    .sout11(sout61_17), .sout12(sout61_18), .sout13(sout61_19), .sout14(sout61_20),
                    .sout21(sout62_17), .sout22(sout62_18), .sout23(sout62_19), .sout24(sout62_20),
                    .sout31(sout63_17), .sout32(sout63_18), .sout33(sout63_19), .sout34(sout63_20),
                    .sout41(sout64_17), .sout42(sout64_18), .sout43(sout64_19), .sout44(sout64_20)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_16_6 (.clk(clk), .rst(rst),
                    .ain1(aout61_20), .ain2(aout62_20), .ain3(aout63_20), .ain4(aout64_20),
                    .win1(wout60_21), .win2(wout60_22), .win3(wout60_23), .win4(wout60_24),
                    .aout1(aout61_24), .aout2(aout62_24), .aout3(aout63_24), .aout4(aout64_24),
                    .wout1(wout64_21), .wout2(wout64_22), .wout3(wout64_23), .wout4(wout64_24),
                    .sout11(sout61_21), .sout12(sout61_22), .sout13(sout61_23), .sout14(sout61_24),
                    .sout21(sout62_21), .sout22(sout62_22), .sout23(sout62_23), .sout24(sout62_24),
                    .sout31(sout63_21), .sout32(sout63_22), .sout33(sout63_23), .sout34(sout63_24),
                    .sout41(sout64_21), .sout42(sout64_22), .sout43(sout64_23), .sout44(sout64_24)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16_7 (.clk(clk), .rst(rst),
                    .ain1(aout61_24), .ain2(aout62_24), .ain3(aout63_24), .ain4(aout64_24),
                    .win1(wout60_25), .win2(wout60_26), .win3(wout60_27), .win4(wout60_28),
                    .aout1(aout61_28), .aout2(aout62_28), .aout3(aout63_28), .aout4(aout64_28),
                    .wout1(wout64_25), .wout2(wout64_26), .wout3(wout64_27), .wout4(wout64_28),
                    .sout11(sout61_25), .sout12(sout61_26), .sout13(sout61_27), .sout14(sout61_28),
                    .sout21(sout62_25), .sout22(sout62_26), .sout23(sout62_27), .sout24(sout62_28),
                    .sout31(sout63_25), .sout32(sout63_26), .sout33(sout63_27), .sout34(sout63_28),
                    .sout41(sout64_25), .sout42(sout64_26), .sout43(sout64_27), .sout44(sout64_28)
                    ); //4x4 MAC array
    
    mac_array_4x4 mac_array_4x4_16_8 (.clk(clk), .rst(rst),
                    .ain1(aout61_28), .ain2(aout62_28), .ain3(aout63_28), .ain4(aout64_28),
                    .win1(wout60_29), .win2(wout60_30), .win3(wout60_31), .win4(wout60_32),
                    .aout1(aout61_32), .aout2(aout62_32), .aout3(aout63_32), .aout4(aout64_32),
                    .wout1(wout64_29), .wout2(wout64_30), .wout3(wout64_31), .wout4(wout64_32),
                    .sout11(sout61_29), .sout12(sout61_30), .sout13(sout61_31), .sout14(sout61_32),
                    .sout21(sout62_29), .sout22(sout62_30), .sout23(sout62_31), .sout24(sout62_32),
                    .sout31(sout63_29), .sout32(sout63_30), .sout33(sout63_31), .sout34(sout63_32),
                    .sout41(sout64_29), .sout42(sout64_30), .sout43(sout64_31), .sout44(sout64_32)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16_9 (.clk(clk), .rst(rst),
                    .ain1(aout61_32), .ain2(aout62_32), .ain3(aout63_32), .ain4(aout64_32),
                    .win1(wout60_33), .win2(wout60_34), .win3(wout60_35), .win4(wout60_36),
                    .aout1(aout61_36), .aout2(aout62_36), .aout3(aout63_36), .aout4(aout64_36),
                    .wout1(wout64_33), .wout2(wout64_34), .wout3(wout64_35), .wout4(wout64_36),
                    .sout11(sout61_33), .sout12(sout61_34), .sout13(sout61_35), .sout14(sout61_36),
                    .sout21(sout62_33), .sout22(sout62_34), .sout23(sout62_35), .sout24(sout62_36),
                    .sout31(sout63_33), .sout32(sout63_34), .sout33(sout63_35), .sout34(sout63_36),
                    .sout41(sout64_33), .sout42(sout64_34), .sout43(sout64_35), .sout44(sout64_36)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16_10 (.clk(clk), .rst(rst),
                    .ain1(aout61_36), .ain2(aout62_36), .ain3(aout63_36), .ain4(aout64_36),
                    .win1(wout60_37), .win2(wout60_38), .win3(wout60_39), .win4(wout60_40),
                    .aout1(aout61_40), .aout2(aout62_40), .aout3(aout63_40), .aout4(aout64_40),
                    .wout1(wout64_37), .wout2(wout64_38), .wout3(wout64_39), .wout4(wout64_40),
                    .sout11(sout61_37), .sout12(sout61_38), .sout13(sout61_39), .sout14(sout61_40),
                    .sout21(sout62_37), .sout22(sout62_38), .sout23(sout62_39), .sout24(sout62_40),
                    .sout31(sout63_37), .sout32(sout63_38), .sout33(sout63_39), .sout34(sout63_40),
                    .sout41(sout64_37), .sout42(sout64_38), .sout43(sout64_39), .sout44(sout64_40)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16_11 (.clk(clk), .rst(rst),
                    .ain1(aout61_40), .ain2(aout62_40), .ain3(aout63_40), .ain4(aout64_40),
                    .win1(wout60_41), .win2(wout60_42), .win3(wout60_43), .win4(wout60_44),
                    .aout1(aout61_44), .aout2(aout62_44), .aout3(aout63_44), .aout4(aout64_44),
                    .wout1(wout64_41), .wout2(wout64_42), .wout3(wout64_43), .wout4(wout64_44),
                    .sout11(sout61_41), .sout12(sout61_42), .sout13(sout61_43), .sout14(sout61_44),
                    .sout21(sout62_41), .sout22(sout62_42), .sout23(sout62_43), .sout24(sout62_44),
                    .sout31(sout63_41), .sout32(sout63_42), .sout33(sout63_43), .sout34(sout63_44),
                    .sout41(sout64_41), .sout42(sout64_42), .sout43(sout64_43), .sout44(sout64_44)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16_12 (.clk(clk), .rst(rst),
                    .ain1(aout61_44), .ain2(aout62_44), .ain3(aout63_44), .ain4(aout64_44),
                    .win1(wout60_45), .win2(wout60_46), .win3(wout60_47), .win4(wout60_48),
                    .aout1(aout61_48), .aout2(aout62_48), .aout3(aout63_48), .aout4(aout64_48),
                    .wout1(wout64_45), .wout2(wout64_46), .wout3(wout64_47), .wout4(wout64_48),
                    .sout11(sout61_45), .sout12(sout61_46), .sout13(sout61_47), .sout14(sout61_48),
                    .sout21(sout62_45), .sout22(sout62_46), .sout23(sout62_47), .sout24(sout62_48),
                    .sout31(sout63_45), .sout32(sout63_46), .sout33(sout63_47), .sout34(sout63_48),
                    .sout41(sout64_45), .sout42(sout64_46), .sout43(sout64_47), .sout44(sout64_48)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16_13 (.clk(clk), .rst(rst),
                    .ain1(aout61_48), .ain2(aout62_48), .ain3(aout63_48), .ain4(aout64_48),
                    .win1(wout60_49), .win2(wout60_50), .win3(wout60_51), .win4(wout60_52),
                    .aout1(aout61_52), .aout2(aout62_52), .aout3(aout63_52), .aout4(aout64_52),
                    .wout1(wout64_49), .wout2(wout64_50), .wout3(wout64_51), .wout4(wout64_52),
                    .sout11(sout61_49), .sout12(sout61_50), .sout13(sout61_51), .sout14(sout61_52),
                    .sout21(sout62_49), .sout22(sout62_50), .sout23(sout62_51), .sout24(sout62_52),
                    .sout31(sout63_49), .sout32(sout63_50), .sout33(sout63_51), .sout34(sout63_52),
                    .sout41(sout64_49), .sout42(sout64_50), .sout43(sout64_51), .sout44(sout64_52)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16_14 (.clk(clk), .rst(rst),
                    .ain1(aout61_52), .ain2(aout62_52), .ain3(aout63_52), .ain4(aout64_52),
                    .win1(wout60_53), .win2(wout60_54), .win3(wout60_55), .win4(wout60_56),
                    .aout1(aout61_56), .aout2(aout62_56), .aout3(aout63_56), .aout4(aout64_56),
                    .wout1(wout64_53), .wout2(wout64_54), .wout3(wout64_55), .wout4(wout64_56),
                    .sout11(sout61_53), .sout12(sout61_54), .sout13(sout61_55), .sout14(sout61_56),
                    .sout21(sout62_53), .sout22(sout62_54), .sout23(sout62_55), .sout24(sout62_56),
                    .sout31(sout63_53), .sout32(sout63_54), .sout33(sout63_55), .sout34(sout63_56),
                    .sout41(sout64_53), .sout42(sout64_54), .sout43(sout64_55), .sout44(sout64_56)
                    ); //4x4 MAC array
                   
    mac_array_4x4 mac_array_4x4_16_15 (.clk(clk), .rst(rst),
                    .ain1(aout61_56), .ain2(aout62_56), .ain3(aout63_56), .ain4(aout64_56),
                    .win1(wout60_57), .win2(wout60_58), .win3(wout60_59), .win4(wout60_60),
                    .aout1(aout61_60), .aout2(aout62_60), .aout3(aout63_60), .aout4(aout64_60),
                    .wout1(wout64_57), .wout2(wout64_58), .wout3(wout64_59), .wout4(wout64_60),
                    .sout11(sout61_57), .sout12(sout61_58), .sout13(sout61_59), .sout14(sout61_60),
                    .sout21(sout62_57), .sout22(sout62_58), .sout23(sout62_59), .sout24(sout62_60),
                    .sout31(sout63_57), .sout32(sout63_58), .sout33(sout63_59), .sout34(sout63_60),
                    .sout41(sout64_57), .sout42(sout64_58), .sout43(sout64_59), .sout44(sout64_60)
                    ); //4x4 MAC array
                    
    mac_array_4x4 mac_array_4x4_16_16 (.clk(clk), .rst(rst),
                    .ain1(aout61_60), .ain2(aout62_60), .ain3(aout63_60), .ain4(aout64_60),
                    .win1(wout60_61), .win2(wout60_62), .win3(wout60_63), .win4(wout60_64),
                    .aout1(aout61_64), .aout2(aout62_64), .aout3(aout63_64), .aout4(aout64_64),
                    .wout1(wout64_61), .wout2(wout64_62), .wout3(wout64_63), .wout4(wout64_64),
                    .sout11(sout61_61), .sout12(sout61_62), .sout13(sout61_63), .sout14(sout61_64),
                    .sout21(sout62_61), .sout22(sout62_62), .sout23(sout62_63), .sout24(sout62_64),
                    .sout31(sout63_61), .sout32(sout63_62), .sout33(sout63_63), .sout34(sout63_64),
                    .sout41(sout64_61), .sout42(sout64_62), .sout43(sout64_63), .sout44(sout64_64)
                    ); //4x4 MAC array
    
endmodule
